`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module RetimeWrapper(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out
);
  wire  sr_out;
  wire  sr_in;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF(
  input        clock,
  input        reset,
  input  [6:0] io_input_0_data,
  input        io_input_0_enable,
  input        io_input_0_reset,
  output [6:0] io_output_data
);
  reg [6:0] ff;
  reg [31:0] _RAND_0;
  wire [6:0] _T_7;
  wire [6:0] _T_8;
  wire [6:0] _T_9;
  assign _T_7 = io_input_0_enable ? io_input_0_data : ff;
  assign _T_8 = io_input_0_reset ? 7'h0 : _T_7;
  assign _T_9 = io_input_0_reset ? 7'h0 : ff;
  assign io_output_data = _T_9;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  ff = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 7'h0;
    end else begin
      if (io_input_0_reset) begin
        ff <= 7'h0;
      end else begin
        if (io_input_0_enable) begin
          ff <= io_input_0_data;
        end
      end
    end
  end
endmodule
module SingleCounter(
  input        clock,
  input        reset,
  input  [6:0] io_input_stop,
  input        io_input_reset,
  input        io_input_enable,
  output       io_output_done
);
  wire  FF_clock;
  wire  FF_reset;
  wire [6:0] FF_io_input_0_data;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [6:0] FF_io_output_data;
  wire [6:0] _T_20;
  wire [7:0] _T_22;
  wire [6:0] _T_23;
  wire [6:0] _T_24;
  wire  _T_27;
  wire [6:0] _T_37;
  wire [6:0] _T_39;
  wire [6:0] _T_40;
  wire  _T_52;
  FF FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  assign _T_20 = $signed(FF_io_output_data);
  assign _T_22 = $signed(_T_20) + $signed(7'sh1);
  assign _T_23 = _T_22[6:0];
  assign _T_24 = $signed(_T_23);
  assign _T_27 = $signed(_T_24) >= $signed(io_input_stop);
  assign _T_37 = _T_27 ? $signed(_T_20) : $signed(_T_24);
  assign _T_39 = $unsigned(_T_37);
  assign _T_40 = io_input_reset ? 7'h0 : _T_39;
  assign _T_52 = io_input_enable & _T_27;
  assign io_output_done = _T_52;
  assign FF_io_input_0_data = _T_40;
  assign FF_io_input_0_enable = io_input_enable;
  assign FF_io_input_0_reset = io_input_reset;
  assign FF_clock = clock;
  assign FF_reset = reset;
endmodule
module SRFF_sp(
  input   clock,
  input   reset,
  input   io_input_set,
  input   io_input_reset,
  input   io_input_asyn_reset,
  output  io_output_data
);
  reg  _T_8;
  reg [31:0] _RAND_0;
  wire  _T_12;
  wire  _T_13;
  wire  _T_14;
  wire  _T_16;
  assign _T_12 = io_input_reset ? 1'h0 : _T_8;
  assign _T_13 = io_input_set ? 1'h1 : _T_12;
  assign _T_14 = io_input_asyn_reset ? 1'h0 : _T_13;
  assign _T_16 = io_input_asyn_reset ? 1'h0 : _T_8;
  assign io_output_data = _T_16;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_8 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_8 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_8 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_8 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_8 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module FF_1(
  input         clock,
  input         reset,
  input  [31:0] io_input_0_data,
  input  [31:0] io_input_0_init,
  input         io_input_0_enable,
  input         io_input_0_reset,
  output [31:0] io_output_data
);
  reg [31:0] ff;
  reg [31:0] _RAND_0;
  wire [31:0] _T_7;
  wire [31:0] _T_8;
  wire [31:0] _T_9;
  assign _T_7 = io_input_0_enable ? io_input_0_data : ff;
  assign _T_8 = io_input_0_reset ? io_input_0_init : _T_7;
  assign _T_9 = io_input_0_reset ? io_input_0_init : ff;
  assign io_output_data = _T_9;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= io_input_0_init;
    end else begin
      if (io_input_0_reset) begin
        ff <= io_input_0_init;
      end else begin
        if (io_input_0_enable) begin
          ff <= io_input_0_data;
        end
      end
    end
  end
endmodule
module RetimeWrapper_1(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  output [31:0] io_out
);
  wire [31:0] sr_out;
  wire [31:0] sr_in;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module SingleCounter_1(
  input         clock,
  input         reset,
  input  [31:0] io_input_stop,
  input         io_input_reset,
  input         io_input_enable,
  output        io_output_done
);
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire [31:0] _T_20;
  wire [32:0] _T_22;
  wire [31:0] _T_23;
  wire [31:0] _T_24;
  wire  _T_27;
  wire [31:0] _T_37;
  wire [31:0] _T_39;
  wire [31:0] _T_40;
  wire  _T_52;
  FF_1 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  assign _T_20 = $signed(FF_io_output_data);
  assign _T_22 = $signed(_T_20) + $signed(32'sh1);
  assign _T_23 = _T_22[31:0];
  assign _T_24 = $signed(_T_23);
  assign _T_27 = $signed(_T_24) >= $signed(io_input_stop);
  assign _T_37 = _T_27 ? $signed(32'sh0) : $signed(_T_24);
  assign _T_39 = $unsigned(_T_37);
  assign _T_40 = io_input_reset ? 32'h0 : _T_39;
  assign _T_52 = io_input_enable & _T_27;
  assign io_output_done = _T_52;
  assign FF_io_input_0_data = _T_40;
  assign FF_io_input_0_init = 32'h0;
  assign FF_io_input_0_enable = io_input_enable;
  assign FF_io_input_0_reset = io_input_reset;
  assign FF_clock = clock;
  assign FF_reset = reset;
endmodule
module Seqpipe(
  input   clock,
  input   reset,
  input   io_input_enable,
  input   io_input_stageDone_0,
  input   io_input_stageDone_1,
  input   io_input_rst,
  output  io_output_done,
  output  io_output_stageEnable_0,
  output  io_output_stageEnable_1,
  output  io_output_rst_en
);
  wire  SingleCounter_clock;
  wire  SingleCounter_reset;
  wire [6:0] SingleCounter_io_input_stop;
  wire  SingleCounter_io_input_reset;
  wire  SingleCounter_io_input_enable;
  wire  SingleCounter_io_output_done;
  wire  SRFF_sp_clock;
  wire  SRFF_sp_reset;
  wire  SRFF_sp_io_input_set;
  wire  SRFF_sp_io_input_reset;
  wire  SRFF_sp_io_input_asyn_reset;
  wire  SRFF_sp_io_output_data;
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire [31:0] _T_25;
  wire  _T_27;
  wire  _T_28;
  wire  _T_30;
  wire  _T_31;
  wire [6:0] _T_35;
  wire  FF_1_clock;
  wire  FF_1_reset;
  wire [31:0] FF_1_io_input_0_data;
  wire [31:0] FF_1_io_input_0_init;
  wire  FF_1_io_input_0_enable;
  wire  FF_1_io_input_0_reset;
  wire [31:0] FF_1_io_output_data;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [31:0] RetimeWrapper_io_in;
  wire [31:0] RetimeWrapper_io_out;
  wire [31:0] _T_42;
  wire  SingleCounter_1_clock;
  wire  SingleCounter_1_reset;
  wire [31:0] SingleCounter_1_io_input_stop;
  wire  SingleCounter_1_io_input_reset;
  wire  SingleCounter_1_io_input_enable;
  wire  SingleCounter_1_io_output_done;
  wire  _T_43;
  wire [31:0] _T_45;
  wire  _T_47;
  wire  _T_48;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_53;
  wire [1:0] _T_65;
  wire [2:0] _T_66;
  wire  _T_70;
  wire [32:0] _T_78;
  wire [31:0] _T_79;
  wire [31:0] _T_80;
  wire [31:0] _T_81;
  wire  _T_83;
  wire  _T_84;
  wire  _T_85;
  wire  _T_86;
  wire [32:0] _T_88;
  wire [31:0] _T_89;
  wire [31:0] _T_90;
  wire [31:0] _T_91;
  wire [31:0] _T_92;
  wire [31:0] _GEN_0;
  wire  _T_94;
  wire [2:0] _GEN_1;
  wire [31:0] _GEN_2;
  wire [31:0] _GEN_3;
  wire [31:0] _GEN_4;
  wire [31:0] _GEN_5;
  wire [31:0] _GEN_6;
  wire [31:0] _GEN_8;
  wire  _T_118;
  SingleCounter SingleCounter (
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_stop(SingleCounter_io_input_stop),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_input_enable(SingleCounter_io_input_enable),
    .io_output_done(SingleCounter_io_output_done)
  );
  SRFF_sp SRFF_sp (
    .clock(SRFF_sp_clock),
    .reset(SRFF_sp_reset),
    .io_input_set(SRFF_sp_io_input_set),
    .io_input_reset(SRFF_sp_io_input_reset),
    .io_input_asyn_reset(SRFF_sp_io_input_asyn_reset),
    .io_output_data(SRFF_sp_io_output_data)
  );
  FF_1 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  FF_1 FF_1 (
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_input_0_data(FF_1_io_input_0_data),
    .io_input_0_init(FF_1_io_input_0_init),
    .io_input_0_enable(FF_1_io_input_0_enable),
    .io_input_0_reset(FF_1_io_input_0_reset),
    .io_output_data(FF_1_io_output_data)
  );
  RetimeWrapper_1 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SingleCounter_1 SingleCounter_1 (
    .clock(SingleCounter_1_clock),
    .reset(SingleCounter_1_reset),
    .io_input_stop(SingleCounter_1_io_input_stop),
    .io_input_reset(SingleCounter_1_io_input_reset),
    .io_input_enable(SingleCounter_1_io_input_enable),
    .io_output_done(SingleCounter_1_io_output_done)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_25 = $signed(FF_io_output_data);
  assign _T_27 = $signed(_T_25) == $signed(32'sh1);
  assign _T_28 = _T_27 & io_input_enable;
  assign _T_30 = $signed(_T_25) != $signed(32'sh1);
  assign _T_31 = _T_30 | io_input_rst;
  assign _T_35 = SRFF_sp_io_output_data ? $signed(7'sh1) : $signed(7'sh1c);
  assign _T_43 = io_input_enable & io_input_stageDone_1;
  assign _T_45 = $signed(_T_42);
  assign _T_47 = $signed(_T_25) == $signed(32'sh4);
  assign _T_48 = io_input_rst | _T_47;
  assign _T_65 = SingleCounter_io_output_done ? 2'h2 : 2'h1;
  assign _T_66 = {{1'd0}, _T_65};
  assign _T_70 = $signed(_T_25) < $signed(32'sh3);
  assign _T_78 = $signed(_T_25) - $signed(32'sh2);
  assign _T_79 = _T_78[31:0];
  assign _T_80 = $signed(_T_79);
  assign _T_81 = $unsigned(_T_80);
  assign _T_83 = 32'h1 == _T_81;
  assign _T_84 = _T_83 ? io_input_stageDone_1 : 1'h0;
  assign _T_85 = 32'h0 == _T_81;
  assign _T_86 = _T_85 ? io_input_stageDone_0 : _T_84;
  assign _T_88 = $signed(_T_25) + $signed(32'sh1);
  assign _T_89 = _T_88[31:0];
  assign _T_90 = $signed(_T_89);
  assign _T_91 = $unsigned(_T_90);
  assign _T_92 = $unsigned(_T_25);
  assign _GEN_0 = _T_86 ? _T_91 : _T_92;
  assign _T_94 = $signed(_T_25) == $signed(32'sh3);
  assign _GEN_1 = SingleCounter_1_io_output_done ? 3'h4 : 3'h2;
  assign _GEN_2 = io_input_stageDone_1 ? {{29'd0}, _GEN_1} : _T_92;
  assign _GEN_3 = _T_47 ? 32'h1 : _T_92;
  assign _GEN_4 = _T_94 ? _GEN_2 : _GEN_3;
  assign _GEN_5 = _T_70 ? _GEN_0 : _GEN_4;
  assign _GEN_6 = _T_27 ? {{29'd0}, _T_66} : _GEN_5;
  assign _GEN_8 = io_input_enable ? _GEN_6 : 32'h1;
  assign _T_118 = $signed(_T_25) == $signed(32'sh2);
  assign io_output_done = _T_47;
  assign io_output_stageEnable_0 = _T_118;
  assign io_output_stageEnable_1 = _T_94;
  assign io_output_rst_en = _T_53;
  assign SingleCounter_io_input_stop = _T_35;
  assign SingleCounter_io_input_reset = _T_31;
  assign SingleCounter_io_input_enable = _T_28;
  assign SingleCounter_clock = clock;
  assign SingleCounter_reset = reset;
  assign SRFF_sp_io_input_set = SingleCounter_io_output_done;
  assign SRFF_sp_io_input_reset = reset;
  assign SRFF_sp_io_input_asyn_reset = reset;
  assign SRFF_sp_clock = clock;
  assign SRFF_sp_reset = reset;
  assign FF_io_input_0_data = _GEN_8;
  assign FF_io_input_0_init = 32'h1;
  assign FF_io_input_0_enable = 1'h1;
  assign FF_io_input_0_reset = io_input_rst;
  assign FF_clock = clock;
  assign FF_reset = reset;
  assign FF_1_io_input_0_data = 32'h1;
  assign FF_1_io_input_0_init = 32'h0;
  assign FF_1_io_input_0_enable = io_input_enable;
  assign FF_1_io_input_0_reset = io_input_rst;
  assign FF_1_clock = clock;
  assign FF_1_reset = reset;
  assign RetimeWrapper_io_in = FF_1_io_output_data;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_42 = RetimeWrapper_io_out;
  assign SingleCounter_1_io_input_stop = _T_45;
  assign SingleCounter_1_io_input_reset = _T_48;
  assign SingleCounter_1_io_input_enable = _T_43;
  assign SingleCounter_1_clock = clock;
  assign SingleCounter_1_reset = reset;
  assign RetimeWrapper_1_io_in = _T_27;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_53 = RetimeWrapper_1_io_out;
endmodule
module SingleCounter_2(
  input   clock,
  input   reset,
  input   io_input_reset,
  input   io_input_enable,
  output  io_output_done
);
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire [31:0] _T_20;
  wire [32:0] _T_22;
  wire [31:0] _T_23;
  wire [31:0] _T_24;
  wire  _T_28;
  wire [31:0] _T_39;
  wire [31:0] _T_41;
  wire [31:0] _T_42;
  wire  _T_55;
  FF_1 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  assign _T_20 = $signed(FF_io_output_data);
  assign _T_22 = $signed(_T_20) + $signed(32'sh1);
  assign _T_23 = _T_22[31:0];
  assign _T_24 = $signed(_T_23);
  assign _T_28 = $signed(_T_24) >= $signed(32'sh1);
  assign _T_39 = _T_28 ? $signed(_T_20) : $signed(_T_24);
  assign _T_41 = $unsigned(_T_39);
  assign _T_42 = io_input_reset ? 32'h0 : _T_41;
  assign _T_55 = io_input_enable & _T_28;
  assign io_output_done = _T_55;
  assign FF_io_input_0_data = _T_42;
  assign FF_io_input_0_init = 32'h0;
  assign FF_io_input_0_enable = io_input_enable;
  assign FF_io_input_0_reset = io_input_reset;
  assign FF_clock = clock;
  assign FF_reset = reset;
endmodule
module Innerpipe(
  input   clock,
  input   reset,
  input   io_input_enable,
  input   io_input_ctr_done,
  input   io_input_rst,
  output  io_output_done,
  output  io_output_ctr_inc
);
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire  SingleCounter_clock;
  wire  SingleCounter_reset;
  wire  SingleCounter_io_input_reset;
  wire  SingleCounter_io_input_enable;
  wire  SingleCounter_io_output_done;
  wire  _T_20;
  wire  _T_21;
  wire  _T_23;
  wire  _T_25;
  wire  _T_26;
  wire  _T_27;
  wire [1:0] _T_42;
  wire [1:0] _T_45;
  wire [1:0] _GEN_0;
  wire  _T_47;
  wire  _GEN_3;
  wire  _T_61;
  wire  _T_69;
  wire [32:0] _T_77;
  wire [31:0] _T_78;
  wire [31:0] _T_79;
  wire [31:0] _GEN_9;
  wire  _GEN_10;
  wire  _GEN_11;
  wire [31:0] _GEN_13;
  wire  _GEN_14;
  wire  _GEN_16;
  wire [31:0] _GEN_17;
  wire  _T_82;
  wire  _T_83;
  wire  _GEN_18;
  wire  _GEN_20;
  wire [31:0] _GEN_21;
  FF_1 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  SingleCounter_2 SingleCounter (
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_input_enable(SingleCounter_io_input_enable),
    .io_output_done(SingleCounter_io_output_done)
  );
  assign _T_20 = FF_io_output_data == 32'h1;
  assign _T_21 = _T_20 & io_input_enable;
  assign _T_23 = FF_io_output_data != 32'h1;
  assign _T_25 = FF_io_output_data < 32'h4;
  assign _T_26 = _T_23 & _T_25;
  assign _T_27 = _T_26 | io_input_rst;
  assign _T_42 = io_input_ctr_done ? 2'h3 : 2'h1;
  assign _T_45 = io_input_ctr_done ? 2'h3 : 2'h2;
  assign _GEN_0 = SingleCounter_io_output_done ? _T_45 : _T_42;
  assign _T_47 = FF_io_output_data == 32'h2;
  assign _GEN_3 = io_input_ctr_done ? 1'h0 : 1'h1;
  assign _T_61 = FF_io_output_data == 32'h3;
  assign _T_69 = FF_io_output_data >= 32'h4;
  assign _T_77 = FF_io_output_data + 32'h1;
  assign _T_78 = _T_77[31:0];
  assign _T_79 = _T_69 ? 32'h1 : _T_78;
  assign _GEN_9 = _T_61 ? 32'h1 : _T_79;
  assign _GEN_10 = _T_47 ? _GEN_3 : 1'h0;
  assign _GEN_11 = _T_47 ? io_input_ctr_done : 1'h0;
  assign _GEN_13 = _T_47 ? {{30'd0}, _T_45} : _GEN_9;
  assign _GEN_14 = _T_20 ? 1'h0 : _GEN_11;
  assign _GEN_16 = _T_20 ? 1'h0 : _GEN_10;
  assign _GEN_17 = _T_20 ? {{30'd0}, _GEN_0} : _GEN_13;
  assign _T_82 = _T_47 & io_input_ctr_done;
  assign _T_83 = io_input_ctr_done | _T_82;
  assign _GEN_18 = io_input_enable ? _GEN_14 : _T_83;
  assign _GEN_20 = io_input_enable ? _GEN_16 : 1'h0;
  assign _GEN_21 = io_input_enable ? _GEN_17 : 32'h1;
  assign io_output_done = _GEN_18;
  assign io_output_ctr_inc = _GEN_20;
  assign FF_io_input_0_data = _GEN_21;
  assign FF_io_input_0_init = 32'h1;
  assign FF_io_input_0_enable = 1'h1;
  assign FF_io_input_0_reset = 1'h0;
  assign FF_clock = clock;
  assign FF_reset = reset;
  assign SingleCounter_io_input_reset = _T_27;
  assign SingleCounter_io_input_enable = _T_21;
  assign SingleCounter_clock = clock;
  assign SingleCounter_reset = reset;
endmodule
module SingleCounter_4(
  input   clock,
  input   reset,
  input   io_input_reset,
  output  io_output_done
);
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_input_0_data;
  wire [31:0] FF_io_input_0_init;
  wire  FF_io_input_0_enable;
  wire  FF_io_input_0_reset;
  wire [31:0] FF_io_output_data;
  wire [31:0] _T_20;
  wire [32:0] _T_22;
  wire [31:0] _T_23;
  wire [31:0] _T_24;
  wire  _T_28;
  wire [31:0] _T_39;
  wire [31:0] _T_41;
  wire [31:0] _T_42;
  FF_1 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_input_0_data(FF_io_input_0_data),
    .io_input_0_init(FF_io_input_0_init),
    .io_input_0_enable(FF_io_input_0_enable),
    .io_input_0_reset(FF_io_input_0_reset),
    .io_output_data(FF_io_output_data)
  );
  assign _T_20 = $signed(FF_io_output_data);
  assign _T_22 = $signed(_T_20) + $signed(32'sh1);
  assign _T_23 = _T_22[31:0];
  assign _T_24 = $signed(_T_23);
  assign _T_28 = $signed(_T_24) >= $signed(32'sh0);
  assign _T_39 = _T_28 ? $signed(_T_20) : $signed(_T_24);
  assign _T_41 = $unsigned(_T_39);
  assign _T_42 = io_input_reset ? 32'h0 : _T_41;
  assign io_output_done = _T_28;
  assign FF_io_input_0_data = _T_42;
  assign FF_io_input_0_init = 32'h0;
  assign FF_io_input_0_enable = 1'h1;
  assign FF_io_input_0_reset = io_input_reset;
  assign FF_clock = clock;
  assign FF_reset = reset;
endmodule
module AccelTop(
  input         clock,
  input         reset,
  input         io_enable,
  output        io_done,
  input  [63:0] io_argIns_0,
  output        io_argOuts_0_valid,
  output [63:0] io_argOuts_0_bits
);
  wire [63:0] x323_data_options_0;
  wire  x323_en_options_0;
  wire  RootController_done;
  wire  RootController_en;
  wire  RootController_resetter;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  retime_released;
  wire  x326_done;
  wire  x326_en;
  wire  x326_base_en;
  wire  x326_resetter;
  wire  x330_done;
  wire  x330_en;
  wire  x330_base_en;
  wire  x330_resetter;
  wire  x330_datapath_en;
  wire  x330_ctr_trivial;
  wire [31:0] x327_number;
  wire [31:0] x328_number;
  wire  RootController_sm_clock;
  wire  RootController_sm_reset;
  wire  RootController_sm_io_input_enable;
  wire  RootController_sm_io_input_stageDone_0;
  wire  RootController_sm_io_input_stageDone_1;
  wire  RootController_sm_io_input_rst;
  wire  RootController_sm_io_output_done;
  wire  RootController_sm_io_output_stageEnable_0;
  wire  RootController_sm_io_output_stageEnable_1;
  wire  RootController_sm_io_output_rst_en;
  wire  x326_sm_clock;
  wire  x326_sm_reset;
  wire  x326_sm_io_input_enable;
  wire  x326_sm_io_input_ctr_done;
  wire  x326_sm_io_input_rst;
  wire  x326_sm_io_output_done;
  wire  x326_sm_io_output_ctr_inc;
  wire  x330_sm_clock;
  wire  x330_sm_reset;
  wire  x330_sm_io_input_enable;
  wire  x330_sm_io_input_ctr_done;
  wire  x330_sm_io_input_rst;
  wire  x330_sm_io_output_done;
  wire  x330_sm_io_output_ctr_inc;
  wire  _T_490;
  wire  _T_492;
  wire  _T_501;
  wire  _T_502;
  wire  retime_counter_clock;
  wire  retime_counter_reset;
  wire  retime_counter_io_input_reset;
  wire  retime_counter_io_output_done;
  wire  RetimeWrapper_1_clock;
  wire  RetimeWrapper_1_reset;
  wire  RetimeWrapper_1_io_in;
  wire  RetimeWrapper_1_io_out;
  wire  _T_511;
  wire  done_latch_clock;
  wire  done_latch_reset;
  wire  done_latch_io_input_set;
  wire  done_latch_io_input_reset;
  wire  done_latch_io_input_asyn_reset;
  wire  done_latch_io_output_data;
  wire  _T_512;
  wire  _T_514;
  wire  _T_520;
  reg  _T_523;
  reg [31:0] _RAND_0;
  wire  _T_529;
  reg  _T_532;
  reg [31:0] _RAND_1;
  wire  RetimeWrapper_2_clock;
  wire  RetimeWrapper_2_reset;
  wire  RetimeWrapper_2_io_in;
  wire  RetimeWrapper_2_io_out;
  wire  _T_549;
  wire  _T_551;
  wire  _T_553;
  wire  _T_554;
  wire  _T_555;
  wire  _T_556;
  wire  _T_557;
  reg  _T_560;
  reg [31:0] _RAND_2;
  wire  _T_566;
  reg  _T_569;
  reg [31:0] _RAND_3;
  wire  RetimeWrapper_3_clock;
  wire  RetimeWrapper_3_reset;
  wire  RetimeWrapper_3_io_in;
  wire  RetimeWrapper_3_io_out;
  wire  _T_579;
  wire  _T_581;
  wire  RetimeWrapper_4_clock;
  wire  RetimeWrapper_4_reset;
  wire  RetimeWrapper_4_io_in;
  wire  RetimeWrapper_4_io_out;
  wire  _T_588;
  wire  _T_590;
  wire  RetimeWrapper_5_clock;
  wire  RetimeWrapper_5_reset;
  wire  RetimeWrapper_5_io_in;
  wire  RetimeWrapper_5_io_out;
  wire  _T_593;
  wire  _T_595;
  wire  _T_596;
  wire  _T_597;
  wire  RetimeWrapper_6_clock;
  wire  RetimeWrapper_6_reset;
  wire  RetimeWrapper_6_io_in;
  wire  RetimeWrapper_6_io_out;
  wire  _T_600;
  wire  _T_602;
  wire  RetimeWrapper_7_clock;
  wire  RetimeWrapper_7_reset;
  wire  RetimeWrapper_7_io_in;
  wire  RetimeWrapper_7_io_out;
  wire  _T_605;
  wire  _T_607;
  wire  _T_608;
  wire  _T_609;
  wire [32:0] _T_615_number;
  wire [32:0] _T_617_number;
  wire [32:0] _T_627;
  wire  _T_630;
  wire [32:0] _T_632;
  wire [33:0] _T_646;
  wire [32:0] _T_647;
  wire [31:0] _T_649_number;
  wire [31:0] _T_663;
  wire [31:0] _T_667;
  wire  _T_668;
  wire [31:0] _T_672;
  wire [63:0] _T_673;
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  Seqpipe RootController_sm (
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_input_enable(RootController_sm_io_input_enable),
    .io_input_stageDone_0(RootController_sm_io_input_stageDone_0),
    .io_input_stageDone_1(RootController_sm_io_input_stageDone_1),
    .io_input_rst(RootController_sm_io_input_rst),
    .io_output_done(RootController_sm_io_output_done),
    .io_output_stageEnable_0(RootController_sm_io_output_stageEnable_0),
    .io_output_stageEnable_1(RootController_sm_io_output_stageEnable_1),
    .io_output_rst_en(RootController_sm_io_output_rst_en)
  );
  Innerpipe x326_sm (
    .clock(x326_sm_clock),
    .reset(x326_sm_reset),
    .io_input_enable(x326_sm_io_input_enable),
    .io_input_ctr_done(x326_sm_io_input_ctr_done),
    .io_input_rst(x326_sm_io_input_rst),
    .io_output_done(x326_sm_io_output_done),
    .io_output_ctr_inc(x326_sm_io_output_ctr_inc)
  );
  Innerpipe x330_sm (
    .clock(x330_sm_clock),
    .reset(x330_sm_reset),
    .io_input_enable(x330_sm_io_input_enable),
    .io_input_ctr_done(x330_sm_io_input_ctr_done),
    .io_input_rst(x330_sm_io_input_rst),
    .io_output_done(x330_sm_io_output_done),
    .io_output_ctr_inc(x330_sm_io_output_ctr_inc)
  );
  SingleCounter_4 retime_counter (
    .clock(retime_counter_clock),
    .reset(retime_counter_reset),
    .io_input_reset(retime_counter_io_input_reset),
    .io_output_done(retime_counter_io_output_done)
  );
  RetimeWrapper RetimeWrapper_1 (
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  SRFF_sp done_latch (
    .clock(done_latch_clock),
    .reset(done_latch_reset),
    .io_input_set(done_latch_io_input_set),
    .io_input_reset(done_latch_io_input_reset),
    .io_input_asyn_reset(done_latch_io_input_asyn_reset),
    .io_output_data(done_latch_io_output_data)
  );
  RetimeWrapper RetimeWrapper_2 (
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 (
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 (
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 (
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 (
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 (
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign _T_490 = RootController_en & retime_released;
  assign _T_492 = retime_released ? RootController_sm_io_output_done : 1'h0;
  assign _T_501 = io_done == 1'h0;
  assign _T_502 = io_enable & _T_501;
  assign _T_512 = x326_en & retime_released;
  assign _T_514 = retime_released ? x326_sm_io_output_done : 1'h0;
  assign _T_520 = ~ x326_sm_io_output_ctr_inc;
  assign _T_529 = x326_sm_io_output_ctr_inc & _T_523;
  assign _T_549 = x330_en & retime_released;
  assign _T_551 = retime_released ? x330_sm_io_output_done : 1'h0;
  assign _T_553 = ~ x330_done;
  assign _T_554 = x330_sm_io_output_ctr_inc & _T_553;
  assign _T_555 = ~ x330_ctr_trivial;
  assign _T_556 = _T_554 & _T_555;
  assign _T_557 = ~ x330_sm_io_output_ctr_inc;
  assign _T_566 = x330_sm_io_output_ctr_inc & _T_560;
  assign _T_581 = retime_released ? _T_579 : 1'h0;
  assign _T_590 = retime_released ? _T_588 : 1'h0;
  assign _T_595 = retime_released ? _T_593 : 1'h0;
  assign _T_596 = ~ _T_595;
  assign _T_597 = _T_590 & _T_596;
  assign _T_602 = retime_released ? _T_600 : 1'h0;
  assign _T_607 = retime_released ? _T_605 : 1'h0;
  assign _T_608 = ~ _T_607;
  assign _T_609 = _T_602 & _T_608;
  assign _T_630 = x327_number[31];
  assign _T_632 = {_T_630,x327_number};
  assign _T_646 = _T_617_number + 33'h4;
  assign _T_647 = _T_646[32:0];
  assign _T_667 = _T_615_number[31:0];
  assign _T_668 = x328_number[31];
  assign _T_672 = _T_668 ? 32'hffffffff : 32'h0;
  assign _T_673 = {_T_672,x328_number};
  assign io_done = done_latch_io_output_data;
  assign io_argOuts_0_valid = x323_en_options_0;
  assign io_argOuts_0_bits = x323_data_options_0;
  assign x323_data_options_0 = _T_673;
  assign x323_en_options_0 = x330_datapath_en;
  assign RootController_done = _T_492;
  assign RootController_en = _T_502;
  assign RootController_resetter = reset;
  assign RetimeWrapper_io_in = 1'h0;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign retime_released = _T_511;
  assign x326_done = _T_514;
  assign x326_en = x326_base_en;
  assign x326_base_en = _T_597;
  assign x326_resetter = RootController_sm_io_output_rst_en;
  assign x330_done = _T_551;
  assign x330_en = x330_base_en;
  assign x330_base_en = _T_609;
  assign x330_resetter = RootController_sm_io_output_rst_en;
  assign x330_datapath_en = _T_556;
  assign x330_ctr_trivial = _T_581;
  assign x327_number = io_argIns_0[31:0];
  assign x328_number = _T_649_number;
  assign RootController_sm_io_input_enable = _T_490;
  assign RootController_sm_io_input_stageDone_0 = x326_done;
  assign RootController_sm_io_input_stageDone_1 = x330_done;
  assign RootController_sm_io_input_rst = RootController_resetter;
  assign RootController_sm_clock = clock;
  assign RootController_sm_reset = reset;
  assign x326_sm_io_input_enable = _T_512;
  assign x326_sm_io_input_ctr_done = _T_532;
  assign x326_sm_io_input_rst = x326_resetter;
  assign x326_sm_clock = clock;
  assign x326_sm_reset = reset;
  assign x330_sm_io_input_enable = _T_549;
  assign x330_sm_io_input_ctr_done = _T_569;
  assign x330_sm_io_input_rst = x330_resetter;
  assign x330_sm_clock = clock;
  assign x330_sm_reset = reset;
  assign retime_counter_io_input_reset = reset;
  assign retime_counter_clock = clock;
  assign retime_counter_reset = reset;
  assign RetimeWrapper_1_io_in = retime_counter_io_output_done;
  assign RetimeWrapper_1_clock = clock;
  assign RetimeWrapper_1_reset = reset;
  assign _T_511 = RetimeWrapper_1_io_out;
  assign done_latch_io_input_set = RootController_done;
  assign done_latch_io_input_reset = RootController_resetter;
  assign done_latch_io_input_asyn_reset = RootController_resetter;
  assign done_latch_clock = clock;
  assign done_latch_reset = reset;
  assign RetimeWrapper_2_io_in = 1'h0;
  assign RetimeWrapper_2_clock = clock;
  assign RetimeWrapper_2_reset = reset;
  assign RetimeWrapper_3_io_in = 1'h0;
  assign RetimeWrapper_3_clock = clock;
  assign RetimeWrapper_3_reset = reset;
  assign _T_579 = RetimeWrapper_3_io_out;
  assign RetimeWrapper_4_io_in = RootController_sm_io_output_stageEnable_0;
  assign RetimeWrapper_4_clock = clock;
  assign RetimeWrapper_4_reset = reset;
  assign _T_588 = RetimeWrapper_4_io_out;
  assign RetimeWrapper_5_io_in = x326_done;
  assign RetimeWrapper_5_clock = clock;
  assign RetimeWrapper_5_reset = reset;
  assign _T_593 = RetimeWrapper_5_io_out;
  assign RetimeWrapper_6_io_in = RootController_sm_io_output_stageEnable_1;
  assign RetimeWrapper_6_clock = clock;
  assign RetimeWrapper_6_reset = reset;
  assign _T_600 = RetimeWrapper_6_io_out;
  assign RetimeWrapper_7_io_in = x330_done;
  assign RetimeWrapper_7_clock = clock;
  assign RetimeWrapper_7_reset = reset;
  assign _T_605 = RetimeWrapper_7_io_out;
  assign _T_615_number = _T_647;
  assign _T_617_number = _T_627;
  assign _T_627 = _T_632;
  assign _T_649_number = _T_663;
  assign _T_663 = _T_667;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_523 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_532 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_560 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_569 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_523 <= 1'h0;
    end else begin
      _T_523 <= _T_520;
    end
    if (reset) begin
      _T_532 <= 1'h0;
    end else begin
      _T_532 <= _T_529;
    end
    if (reset) begin
      _T_560 <= 1'h0;
    end else begin
      _T_560 <= _T_557;
    end
    if (reset) begin
      _T_569 <= 1'h0;
    end else begin
      _T_569 <= _T_566;
    end
  end
endmodule
module FF_9(
  input   clock,
  input   reset,
  input   io_in,
  output  io_out,
  input   io_enable
);
  wire  d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire  RetimeWrapper_io_in;
  wire  RetimeWrapper_io_out;
  wire  _T_9;
  wire  _GEN_0;
  wire  _GEN_1;
  RetimeWrapper RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? 1'h0 : _T_9;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_9;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_9 = RetimeWrapper_io_out;
endmodule
module RetimeWrapper_11(
  input        clock,
  input        reset,
  input  [9:0] io_in,
  output [9:0] io_out
);
  wire [9:0] sr_out;
  wire [9:0] sr_in;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(10), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_10(
  input        clock,
  input        reset,
  input  [9:0] io_in,
  output [9:0] io_out,
  input        io_enable
);
  wire [9:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [9:0] RetimeWrapper_io_in;
  wire [9:0] RetimeWrapper_io_out;
  wire [9:0] _T_9;
  wire [9:0] _GEN_0;
  wire [9:0] _GEN_1;
  RetimeWrapper_11 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? 10'h0 : _T_9;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_9;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_9 = RetimeWrapper_io_out;
endmodule
module UpDownCtr(
  input        clock,
  input        reset,
  input  [9:0] io_strideInc,
  input  [9:0] io_strideDec,
  input        io_dec,
  output [9:0] io_out,
  output [9:0] io_nextInc,
  output [9:0] io_nextDec
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [9:0] reg$_io_in;
  wire [9:0] reg$_io_out;
  wire  reg$_io_enable;
  wire [9:0] decval;
  wire [10:0] _T_20;
  wire [10:0] _T_21;
  wire [9:0] incr;
  wire [10:0] _T_22;
  wire [9:0] newval;
  wire [10:0] _T_27;
  wire [9:0] _T_28;
  wire [10:0] _T_29;
  wire [10:0] _T_30;
  wire [9:0] _T_31;
  FF_10 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign decval = io_dec ? io_strideDec : 10'h0;
  assign _T_20 = 10'h0 - decval;
  assign _T_21 = $unsigned(_T_20);
  assign incr = _T_21[9:0];
  assign _T_22 = reg$_io_out + incr;
  assign newval = _T_22[9:0];
  assign _T_27 = reg$_io_out + io_strideInc;
  assign _T_28 = _T_27[9:0];
  assign _T_29 = reg$_io_out - io_strideDec;
  assign _T_30 = $unsigned(_T_29);
  assign _T_31 = _T_30[9:0];
  assign io_out = reg$_io_out;
  assign io_nextInc = _T_28;
  assign io_nextDec = _T_31;
  assign reg$_io_in = newval;
  assign reg$_io_enable = io_dec;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module Counter(
  input        clock,
  input        reset,
  input  [9:0] io_max,
  output [9:0] io_out,
  output [9:0] io_next,
  input        io_enable,
  output       io_done
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [9:0] reg$_io_in;
  wire [9:0] reg$_io_out;
  wire  reg$_io_enable;
  wire [10:0] count;
  wire [11:0] _T_12;
  wire [10:0] newval;
  wire [10:0] _GEN_1;
  wire  isMax;
  wire [10:0] next;
  wire  _T_14;
  FF_10 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out};
  assign _T_12 = count + 11'h1;
  assign newval = _T_12[10:0];
  assign _GEN_1 = {{1'd0}, io_max};
  assign isMax = newval >= _GEN_1;
  assign next = isMax ? 11'h0 : newval;
  assign _T_14 = io_enable & isMax;
  assign io_out = count[9:0];
  assign io_next = next[9:0];
  assign io_done = _T_14;
  assign reg$_io_in = next[9:0];
  assign reg$_io_enable = io_enable;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module Depulser(
  input   clock,
  input   reset,
  input   io_in,
  input   io_rst,
  output  io_out
);
  wire  r_clock;
  wire  r_reset;
  wire  r_io_in;
  wire  r_io_out;
  wire  r_io_enable;
  wire  _T_6;
  wire  _T_8;
  FF_9 r (
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign _T_6 = io_rst ? 1'h0 : io_in;
  assign _T_8 = io_in | io_rst;
  assign io_out = r_io_out;
  assign r_io_in = _T_6;
  assign r_io_enable = _T_8;
  assign r_clock = clock;
  assign r_reset = reset;
endmodule
module CounterCore(
  input        clock,
  input        reset,
  output [9:0] io_out,
  output [9:0] io_next,
  input        io_enable,
  output       io_done,
  input  [9:0] io_config_max
);
  wire  counter_clock;
  wire  counter_reset;
  wire [9:0] counter_io_max;
  wire [9:0] counter_io_out;
  wire [9:0] counter_io_next;
  wire  counter_io_enable;
  wire  counter_io_done;
  wire  depulser_clock;
  wire  depulser_reset;
  wire  depulser_io_in;
  wire  depulser_io_rst;
  wire  depulser_io_out;
  Counter counter (
    .clock(counter_clock),
    .reset(counter_reset),
    .io_max(counter_io_max),
    .io_out(counter_io_out),
    .io_next(counter_io_next),
    .io_enable(counter_io_enable),
    .io_done(counter_io_done)
  );
  Depulser depulser (
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign io_out = counter_io_out;
  assign io_next = counter_io_next;
  assign io_done = counter_io_done;
  assign counter_io_max = io_config_max;
  assign counter_io_enable = io_enable;
  assign counter_clock = clock;
  assign counter_reset = reset;
  assign depulser_io_in = counter_io_done;
  assign depulser_io_rst = 1'h0;
  assign depulser_clock = clock;
  assign depulser_reset = reset;
endmodule
module CounterChainCore(
  input        clock,
  input        reset,
  output [9:0] io_out_1,
  output [9:0] io_next_1,
  input        io_enable_0,
  output       io_done_0
);
  wire  counters_0_clock;
  wire  counters_0_reset;
  wire [9:0] counters_0_io_out;
  wire [9:0] counters_0_io_next;
  wire  counters_0_io_enable;
  wire  counters_0_io_done;
  wire [9:0] counters_0_io_config_max;
  wire  counters_1_clock;
  wire  counters_1_reset;
  wire [9:0] counters_1_io_out;
  wire [9:0] counters_1_io_next;
  wire  counters_1_io_enable;
  wire  counters_1_io_done;
  wire [9:0] counters_1_io_config_max;
  wire  _T_69;
  CounterCore counters_0 (
    .clock(counters_0_clock),
    .reset(counters_0_reset),
    .io_out(counters_0_io_out),
    .io_next(counters_0_io_next),
    .io_enable(counters_0_io_enable),
    .io_done(counters_0_io_done),
    .io_config_max(counters_0_io_config_max)
  );
  CounterCore counters_1 (
    .clock(counters_1_clock),
    .reset(counters_1_reset),
    .io_out(counters_1_io_out),
    .io_next(counters_1_io_next),
    .io_enable(counters_1_io_enable),
    .io_done(counters_1_io_done),
    .io_config_max(counters_1_io_config_max)
  );
  assign _T_69 = counters_0_io_done;
  assign io_out_1 = counters_1_io_out;
  assign io_next_1 = counters_1_io_next;
  assign io_done_0 = counters_0_io_done;
  assign counters_0_io_enable = io_enable_0;
  assign counters_0_io_config_max = 10'h1;
  assign counters_0_clock = clock;
  assign counters_0_reset = reset;
  assign counters_1_io_enable = _T_69;
  assign counters_1_io_config_max = 10'h200;
  assign counters_1_clock = clock;
  assign counters_1_reset = reset;
endmodule
module SRAM(
  input         clock,
  input  [8:0]  io_raddr,
  input  [8:0]  io_waddr,
  output [81:0] io_rdata
);
  wire [81:0] SRAMVerilogAWS_rdata;
  wire [81:0] SRAMVerilogAWS_wdata;
  wire  SRAMVerilogAWS_wen;
  wire  SRAMVerilogAWS_waddrEn;
  wire  SRAMVerilogAWS_raddrEn;
  wire [8:0] SRAMVerilogAWS_waddr;
  wire [8:0] SRAMVerilogAWS_raddr;
  wire  SRAMVerilogAWS_clk;
  wire [81:0] _T_17;
  SRAMVerilogAWS #(.DWIDTH(82), .WORDS(512), .AWIDTH(9)) SRAMVerilogAWS (
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = SRAMVerilogAWS_rdata;
  assign io_rdata = _T_17;
  assign SRAMVerilogAWS_wdata = 82'h0;
  assign SRAMVerilogAWS_wen = 1'h0;
  assign SRAMVerilogAWS_waddrEn = 1'h1;
  assign SRAMVerilogAWS_raddrEn = 1'h1;
  assign SRAMVerilogAWS_waddr = io_waddr;
  assign SRAMVerilogAWS_raddr = io_raddr;
  assign SRAMVerilogAWS_clk = clock;
endmodule
module MuxN(
  input  [81:0] io_ins_0,
  output [81:0] io_out
);
  assign io_out = io_ins_0;
endmodule
module FIFOCore(
  input         clock,
  input         reset,
  output [81:0] io_deq_0,
  input         io_deqVld,
  output        io_empty,
  output        io_almostEmpty
);
  wire  sizeUDC_clock;
  wire  sizeUDC_reset;
  wire [9:0] sizeUDC_io_strideInc;
  wire [9:0] sizeUDC_io_strideDec;
  wire  sizeUDC_io_dec;
  wire [9:0] sizeUDC_io_out;
  wire [9:0] sizeUDC_io_nextInc;
  wire [9:0] sizeUDC_io_nextDec;
  wire  empty;
  wire  almostEmpty;
  wire  _T_37;
  wire  readEn;
  wire  wptr_clock;
  wire  wptr_reset;
  wire [9:0] wptr_io_out_1;
  wire [9:0] wptr_io_next_1;
  wire  wptr_io_enable_0;
  wire  wptr_io_done_0;
  wire  rptr_clock;
  wire  rptr_reset;
  wire [9:0] rptr_io_out_1;
  wire [9:0] rptr_io_next_1;
  wire  rptr_io_enable_0;
  wire  rptr_io_done_0;
  wire [9:0] nextHeadLocalAddr;
  wire  mems_0_clock;
  wire [8:0] mems_0_io_raddr;
  wire [8:0] mems_0_io_waddr;
  wire [81:0] mems_0_io_rdata;
  wire [9:0] _T_75;
  wire [81:0] MuxN_io_ins_0;
  wire [81:0] MuxN_io_out;
  wire [81:0] _T_84_0;
  UpDownCtr sizeUDC (
    .clock(sizeUDC_clock),
    .reset(sizeUDC_reset),
    .io_strideInc(sizeUDC_io_strideInc),
    .io_strideDec(sizeUDC_io_strideDec),
    .io_dec(sizeUDC_io_dec),
    .io_out(sizeUDC_io_out),
    .io_nextInc(sizeUDC_io_nextInc),
    .io_nextDec(sizeUDC_io_nextDec)
  );
  CounterChainCore wptr (
    .clock(wptr_clock),
    .reset(wptr_reset),
    .io_out_1(wptr_io_out_1),
    .io_next_1(wptr_io_next_1),
    .io_enable_0(wptr_io_enable_0),
    .io_done_0(wptr_io_done_0)
  );
  CounterChainCore rptr (
    .clock(rptr_clock),
    .reset(rptr_reset),
    .io_out_1(rptr_io_out_1),
    .io_next_1(rptr_io_next_1),
    .io_enable_0(rptr_io_enable_0),
    .io_done_0(rptr_io_done_0)
  );
  SRAM mems_0 (
    .clock(mems_0_clock),
    .io_raddr(mems_0_io_raddr),
    .io_waddr(mems_0_io_waddr),
    .io_rdata(mems_0_io_rdata)
  );
  MuxN MuxN (
    .io_ins_0(MuxN_io_ins_0),
    .io_out(MuxN_io_out)
  );
  assign empty = sizeUDC_io_out < 10'h1;
  assign almostEmpty = sizeUDC_io_nextDec < 10'h1;
  assign _T_37 = ~ empty;
  assign readEn = io_deqVld & _T_37;
  assign nextHeadLocalAddr = rptr_io_done_0 ? rptr_io_next_1 : rptr_io_out_1;
  assign _T_75 = readEn ? nextHeadLocalAddr : rptr_io_out_1;
  assign io_deq_0 = MuxN_io_out;
  assign io_empty = empty;
  assign io_almostEmpty = almostEmpty;
  assign sizeUDC_io_strideInc = 10'h1;
  assign sizeUDC_io_strideDec = 10'h1;
  assign sizeUDC_io_dec = readEn;
  assign sizeUDC_clock = clock;
  assign sizeUDC_reset = reset;
  assign wptr_io_enable_0 = 1'h0;
  assign wptr_clock = clock;
  assign wptr_reset = reset;
  assign rptr_io_enable_0 = readEn;
  assign rptr_clock = clock;
  assign rptr_reset = reset;
  assign mems_0_io_raddr = _T_75[8:0];
  assign mems_0_io_waddr = wptr_io_out_1[8:0];
  assign mems_0_clock = clock;
  assign MuxN_io_ins_0 = _T_84_0;
  assign _T_84_0 = mems_0_io_rdata;
endmodule
module MuxVec(
  input  [81:0] io_ins_0_0,
  input  [81:0] io_ins_1_0,
  input         io_sel,
  output [81:0] io_out_0
);
  wire [81:0] _GEN_0_0;
  wire [81:0] _GEN_1;
  assign _GEN_1 = io_sel ? io_ins_1_0 : io_ins_0_0;
  assign io_out_0 = _GEN_0_0;
  assign _GEN_0_0 = _GEN_1;
endmodule
module FIFOArbiter(
  input         clock,
  input         reset,
  output [81:0] io_deq_0,
  input         io_deqVld,
  output        io_empty,
  output        io_tag
);
  wire  tagFF_clock;
  wire  tagFF_reset;
  wire  tagFF_io_in;
  wire  tagFF_io_out;
  wire  tagFF_io_enable;
  wire  tag;
  wire  FIFOCore_clock;
  wire  FIFOCore_reset;
  wire [81:0] FIFOCore_io_deq_0;
  wire  FIFOCore_io_deqVld;
  wire  FIFOCore_io_empty;
  wire  FIFOCore_io_almostEmpty;
  wire  _T_81;
  wire  _T_82;
  wire  FIFOCore_1_clock;
  wire  FIFOCore_1_reset;
  wire [81:0] FIFOCore_1_io_deq_0;
  wire  FIFOCore_1_io_deqVld;
  wire  FIFOCore_1_io_empty;
  wire  FIFOCore_1_io_almostEmpty;
  wire  _T_87;
  wire  _T_89;
  wire  _T_93;
  wire  _T_96;
  wire  _T_99;
  wire  _T_100;
  wire  _T_101;
  wire  _T_114_0;
  wire  _T_119_0;
  wire  _T_129;
  wire [81:0] MuxVec_io_ins_0_0;
  wire [81:0] MuxVec_io_ins_1_0;
  wire  MuxVec_io_sel;
  wire [81:0] MuxVec_io_out_0;
  wire [81:0] _T_147_0_0;
  wire [81:0] _T_147_1_0;
  wire  _T_199;
  wire  _T_200;
  wire  _T_201;
  FF_9 tagFF (
    .clock(tagFF_clock),
    .reset(tagFF_reset),
    .io_in(tagFF_io_in),
    .io_out(tagFF_io_out),
    .io_enable(tagFF_io_enable)
  );
  FIFOCore FIFOCore (
    .clock(FIFOCore_clock),
    .reset(FIFOCore_reset),
    .io_deq_0(FIFOCore_io_deq_0),
    .io_deqVld(FIFOCore_io_deqVld),
    .io_empty(FIFOCore_io_empty),
    .io_almostEmpty(FIFOCore_io_almostEmpty)
  );
  FIFOCore FIFOCore_1 (
    .clock(FIFOCore_1_clock),
    .reset(FIFOCore_1_reset),
    .io_deq_0(FIFOCore_1_io_deq_0),
    .io_deqVld(FIFOCore_1_io_deqVld),
    .io_empty(FIFOCore_1_io_empty),
    .io_almostEmpty(FIFOCore_1_io_almostEmpty)
  );
  MuxVec MuxVec (
    .io_ins_0_0(MuxVec_io_ins_0_0),
    .io_ins_1_0(MuxVec_io_ins_1_0),
    .io_sel(MuxVec_io_sel),
    .io_out_0(MuxVec_io_out_0)
  );
  assign tag = tagFF_io_out;
  assign _T_81 = tag == 1'h0;
  assign _T_82 = io_deqVld & _T_81;
  assign _T_87 = io_deqVld & tag;
  assign _T_89 = FIFOCore_io_empty & FIFOCore_1_io_empty;
  assign _T_93 = FIFOCore_io_empty;
  assign _T_96 = _T_81 & io_deqVld;
  assign _T_99 = _T_96 & FIFOCore_io_almostEmpty;
  assign _T_100 = _T_93 | _T_99;
  assign _T_101 = ~ _T_100;
  assign _T_119_0 = _T_89 ? 1'h0 : _T_114_0;
  assign _T_129 = _T_119_0 ? 1'h0 : 1'h1;
  assign _T_199 = tag ? FIFOCore_1_io_empty : 1'h0;
  assign _T_200 = 1'h0 == tag;
  assign _T_201 = _T_200 ? FIFOCore_io_empty : _T_199;
  assign io_deq_0 = MuxVec_io_out_0;
  assign io_empty = _T_201;
  assign io_tag = tag;
  assign tagFF_io_in = _T_129;
  assign tagFF_io_enable = io_deqVld;
  assign tagFF_clock = clock;
  assign tagFF_reset = reset;
  assign FIFOCore_io_deqVld = _T_82;
  assign FIFOCore_clock = clock;
  assign FIFOCore_reset = reset;
  assign FIFOCore_1_io_deqVld = _T_87;
  assign FIFOCore_1_clock = clock;
  assign FIFOCore_1_reset = reset;
  assign _T_114_0 = _T_101;
  assign MuxVec_io_ins_0_0 = _T_147_0_0;
  assign MuxVec_io_ins_1_0 = _T_147_1_0;
  assign MuxVec_io_sel = tag;
  assign _T_147_0_0 = FIFOCore_io_deq_0;
  assign _T_147_1_0 = FIFOCore_1_io_deq_0;
endmodule
module RetimeWrapper_31(
  input        clock,
  input        reset,
  input  [5:0] io_in,
  output [5:0] io_out
);
  wire [5:0] sr_out;
  wire [5:0] sr_in;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(6), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_32(
  input        clock,
  input        reset,
  output [5:0] io_out
);
  wire [5:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [5:0] RetimeWrapper_io_in;
  wire [5:0] RetimeWrapper_io_out;
  wire [5:0] _T_9;
  wire [5:0] _GEN_0;
  RetimeWrapper_31 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? 6'h0 : _T_9;
  assign io_out = _T_9;
  assign d = _GEN_0;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_9 = RetimeWrapper_io_out;
endmodule
module Counter_8(
  input        clock,
  input        reset,
  output [5:0] io_out
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [5:0] reg$_io_out;
  wire [6:0] count;
  FF_32 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_out(reg$_io_out)
  );
  assign count = {1'h0,reg$_io_out};
  assign io_out = count[5:0];
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module CounterCore_8(
  input        clock,
  input        reset,
  output [5:0] io_out
);
  wire  counter_clock;
  wire  counter_reset;
  wire [5:0] counter_io_out;
  wire  depulser_clock;
  wire  depulser_reset;
  wire  depulser_io_in;
  wire  depulser_io_rst;
  wire  depulser_io_out;
  Counter_8 counter (
    .clock(counter_clock),
    .reset(counter_reset),
    .io_out(counter_io_out)
  );
  Depulser depulser (
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign io_out = counter_io_out;
  assign counter_clock = clock;
  assign counter_reset = reset;
  assign depulser_io_in = 1'h0;
  assign depulser_io_rst = 1'h0;
  assign depulser_clock = clock;
  assign depulser_reset = reset;
endmodule
module CounterChainCore_4(
  input        clock,
  input        reset,
  output [5:0] io_out_0,
  output [5:0] io_out_1
);
  wire  counters_0_clock;
  wire  counters_0_reset;
  wire [5:0] counters_0_io_out;
  wire  counters_1_clock;
  wire  counters_1_reset;
  wire [5:0] counters_1_io_out;
  CounterCore_8 counters_0 (
    .clock(counters_0_clock),
    .reset(counters_0_reset),
    .io_out(counters_0_io_out)
  );
  CounterCore_8 counters_1 (
    .clock(counters_1_clock),
    .reset(counters_1_reset),
    .io_out(counters_1_io_out)
  );
  assign io_out_0 = counters_0_io_out;
  assign io_out_1 = counters_1_io_out;
  assign counters_0_clock = clock;
  assign counters_0_reset = reset;
  assign counters_1_clock = clock;
  assign counters_1_reset = reset;
endmodule
module SRAM_2(
  input        clock,
  input  [4:0] io_raddr,
  input  [4:0] io_waddr
);
  wire [31:0] SRAMVerilogAWS_rdata;
  wire [31:0] SRAMVerilogAWS_wdata;
  wire  SRAMVerilogAWS_wen;
  wire  SRAMVerilogAWS_waddrEn;
  wire  SRAMVerilogAWS_raddrEn;
  wire [4:0] SRAMVerilogAWS_waddr;
  wire [4:0] SRAMVerilogAWS_raddr;
  wire  SRAMVerilogAWS_clk;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(32), .AWIDTH(5)) SRAMVerilogAWS (
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign SRAMVerilogAWS_wdata = 32'h0;
  assign SRAMVerilogAWS_wen = 1'h0;
  assign SRAMVerilogAWS_waddrEn = 1'h1;
  assign SRAMVerilogAWS_raddrEn = 1'h1;
  assign SRAMVerilogAWS_waddr = io_waddr;
  assign SRAMVerilogAWS_raddr = io_raddr;
  assign SRAMVerilogAWS_clk = clock;
endmodule
module RetimeWrapper_39(
  input        clock,
  input        reset,
  input  [3:0] io_in
);
  wire [3:0] sr_out;
  wire [3:0] sr_in;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(4), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign sr_in = io_in;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_40(
  input        clock,
  input        reset,
  input  [3:0] io_in
);
  wire [3:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [3:0] RetimeWrapper_io_in;
  RetimeWrapper_39 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in)
  );
  assign d = io_in;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
endmodule
module FIFOCore_2(
  input   clock,
  input   reset,
  output  io_full,
  output  io_empty,
  output  io_almostFull
);
  wire  sizeUDC_clock;
  wire  sizeUDC_reset;
  wire [9:0] sizeUDC_io_strideInc;
  wire [9:0] sizeUDC_io_strideDec;
  wire  sizeUDC_io_dec;
  wire [9:0] sizeUDC_io_out;
  wire [9:0] sizeUDC_io_nextInc;
  wire [9:0] sizeUDC_io_nextDec;
  wire [10:0] _T_53;
  wire [10:0] _T_54;
  wire [9:0] remainingSlots;
  wire [10:0] _T_56;
  wire [10:0] _T_57;
  wire [9:0] nextRemainingSlots;
  wire  empty;
  wire  full;
  wire  almostFull;
  wire  wptr_clock;
  wire  wptr_reset;
  wire [5:0] wptr_io_out_0;
  wire [5:0] wptr_io_out_1;
  wire  rptr_clock;
  wire  rptr_reset;
  wire [5:0] rptr_io_out_0;
  wire [5:0] rptr_io_out_1;
  wire [5:0] _T_104;
  wire  mems_0_clock;
  wire [4:0] mems_0_io_raddr;
  wire [4:0] mems_0_io_waddr;
  wire  mems_1_clock;
  wire [4:0] mems_1_io_raddr;
  wire [4:0] mems_1_io_waddr;
  wire  mems_2_clock;
  wire [4:0] mems_2_io_raddr;
  wire [4:0] mems_2_io_waddr;
  wire  mems_3_clock;
  wire [4:0] mems_3_io_raddr;
  wire [4:0] mems_3_io_waddr;
  wire  mems_4_clock;
  wire [4:0] mems_4_io_raddr;
  wire [4:0] mems_4_io_waddr;
  wire  mems_5_clock;
  wire [4:0] mems_5_io_raddr;
  wire [4:0] mems_5_io_waddr;
  wire  mems_6_clock;
  wire [4:0] mems_6_io_raddr;
  wire [4:0] mems_6_io_waddr;
  wire  mems_7_clock;
  wire [4:0] mems_7_io_raddr;
  wire [4:0] mems_7_io_waddr;
  wire  mems_8_clock;
  wire [4:0] mems_8_io_raddr;
  wire [4:0] mems_8_io_waddr;
  wire  mems_9_clock;
  wire [4:0] mems_9_io_raddr;
  wire [4:0] mems_9_io_waddr;
  wire  mems_10_clock;
  wire [4:0] mems_10_io_raddr;
  wire [4:0] mems_10_io_waddr;
  wire  mems_11_clock;
  wire [4:0] mems_11_io_raddr;
  wire [4:0] mems_11_io_waddr;
  wire  mems_12_clock;
  wire [4:0] mems_12_io_raddr;
  wire [4:0] mems_12_io_waddr;
  wire  mems_13_clock;
  wire [4:0] mems_13_io_raddr;
  wire [4:0] mems_13_io_waddr;
  wire  mems_14_clock;
  wire [4:0] mems_14_io_raddr;
  wire [4:0] mems_14_io_waddr;
  wire  mems_15_clock;
  wire [4:0] mems_15_io_raddr;
  wire [4:0] mems_15_io_waddr;
  wire  FF_clock;
  wire  FF_reset;
  wire [3:0] FF_io_in;
  wire [5:0] _T_110;
  UpDownCtr sizeUDC (
    .clock(sizeUDC_clock),
    .reset(sizeUDC_reset),
    .io_strideInc(sizeUDC_io_strideInc),
    .io_strideDec(sizeUDC_io_strideDec),
    .io_dec(sizeUDC_io_dec),
    .io_out(sizeUDC_io_out),
    .io_nextInc(sizeUDC_io_nextInc),
    .io_nextDec(sizeUDC_io_nextDec)
  );
  CounterChainCore_4 wptr (
    .clock(wptr_clock),
    .reset(wptr_reset),
    .io_out_0(wptr_io_out_0),
    .io_out_1(wptr_io_out_1)
  );
  CounterChainCore_4 rptr (
    .clock(rptr_clock),
    .reset(rptr_reset),
    .io_out_0(rptr_io_out_0),
    .io_out_1(rptr_io_out_1)
  );
  SRAM_2 mems_0 (
    .clock(mems_0_clock),
    .io_raddr(mems_0_io_raddr),
    .io_waddr(mems_0_io_waddr)
  );
  SRAM_2 mems_1 (
    .clock(mems_1_clock),
    .io_raddr(mems_1_io_raddr),
    .io_waddr(mems_1_io_waddr)
  );
  SRAM_2 mems_2 (
    .clock(mems_2_clock),
    .io_raddr(mems_2_io_raddr),
    .io_waddr(mems_2_io_waddr)
  );
  SRAM_2 mems_3 (
    .clock(mems_3_clock),
    .io_raddr(mems_3_io_raddr),
    .io_waddr(mems_3_io_waddr)
  );
  SRAM_2 mems_4 (
    .clock(mems_4_clock),
    .io_raddr(mems_4_io_raddr),
    .io_waddr(mems_4_io_waddr)
  );
  SRAM_2 mems_5 (
    .clock(mems_5_clock),
    .io_raddr(mems_5_io_raddr),
    .io_waddr(mems_5_io_waddr)
  );
  SRAM_2 mems_6 (
    .clock(mems_6_clock),
    .io_raddr(mems_6_io_raddr),
    .io_waddr(mems_6_io_waddr)
  );
  SRAM_2 mems_7 (
    .clock(mems_7_clock),
    .io_raddr(mems_7_io_raddr),
    .io_waddr(mems_7_io_waddr)
  );
  SRAM_2 mems_8 (
    .clock(mems_8_clock),
    .io_raddr(mems_8_io_raddr),
    .io_waddr(mems_8_io_waddr)
  );
  SRAM_2 mems_9 (
    .clock(mems_9_clock),
    .io_raddr(mems_9_io_raddr),
    .io_waddr(mems_9_io_waddr)
  );
  SRAM_2 mems_10 (
    .clock(mems_10_clock),
    .io_raddr(mems_10_io_raddr),
    .io_waddr(mems_10_io_waddr)
  );
  SRAM_2 mems_11 (
    .clock(mems_11_clock),
    .io_raddr(mems_11_io_raddr),
    .io_waddr(mems_11_io_waddr)
  );
  SRAM_2 mems_12 (
    .clock(mems_12_clock),
    .io_raddr(mems_12_io_raddr),
    .io_waddr(mems_12_io_waddr)
  );
  SRAM_2 mems_13 (
    .clock(mems_13_clock),
    .io_raddr(mems_13_io_raddr),
    .io_waddr(mems_13_io_waddr)
  );
  SRAM_2 mems_14 (
    .clock(mems_14_clock),
    .io_raddr(mems_14_io_raddr),
    .io_waddr(mems_14_io_waddr)
  );
  SRAM_2 mems_15 (
    .clock(mems_15_clock),
    .io_raddr(mems_15_io_raddr),
    .io_waddr(mems_15_io_waddr)
  );
  FF_40 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_in(FF_io_in)
  );
  assign _T_53 = 10'h200 - sizeUDC_io_out;
  assign _T_54 = $unsigned(_T_53);
  assign remainingSlots = _T_54[9:0];
  assign _T_56 = 10'h200 - sizeUDC_io_nextInc;
  assign _T_57 = $unsigned(_T_56);
  assign nextRemainingSlots = _T_57[9:0];
  assign empty = sizeUDC_io_out < 10'h10;
  assign full = remainingSlots < 10'h10;
  assign almostFull = nextRemainingSlots < 10'h10;
  assign _T_104 = rptr_io_out_1;
  assign _T_110 = rptr_io_out_0;
  assign io_full = full;
  assign io_empty = empty;
  assign io_almostFull = almostFull;
  assign sizeUDC_io_strideInc = 10'h10;
  assign sizeUDC_io_strideDec = 10'h10;
  assign sizeUDC_io_dec = 1'h0;
  assign sizeUDC_clock = clock;
  assign sizeUDC_reset = reset;
  assign wptr_clock = clock;
  assign wptr_reset = reset;
  assign rptr_clock = clock;
  assign rptr_reset = reset;
  assign mems_0_io_raddr = _T_104[4:0];
  assign mems_0_io_waddr = wptr_io_out_1[4:0];
  assign mems_0_clock = clock;
  assign mems_1_io_raddr = _T_104[4:0];
  assign mems_1_io_waddr = wptr_io_out_1[4:0];
  assign mems_1_clock = clock;
  assign mems_2_io_raddr = _T_104[4:0];
  assign mems_2_io_waddr = wptr_io_out_1[4:0];
  assign mems_2_clock = clock;
  assign mems_3_io_raddr = _T_104[4:0];
  assign mems_3_io_waddr = wptr_io_out_1[4:0];
  assign mems_3_clock = clock;
  assign mems_4_io_raddr = _T_104[4:0];
  assign mems_4_io_waddr = wptr_io_out_1[4:0];
  assign mems_4_clock = clock;
  assign mems_5_io_raddr = _T_104[4:0];
  assign mems_5_io_waddr = wptr_io_out_1[4:0];
  assign mems_5_clock = clock;
  assign mems_6_io_raddr = _T_104[4:0];
  assign mems_6_io_waddr = wptr_io_out_1[4:0];
  assign mems_6_clock = clock;
  assign mems_7_io_raddr = _T_104[4:0];
  assign mems_7_io_waddr = wptr_io_out_1[4:0];
  assign mems_7_clock = clock;
  assign mems_8_io_raddr = _T_104[4:0];
  assign mems_8_io_waddr = wptr_io_out_1[4:0];
  assign mems_8_clock = clock;
  assign mems_9_io_raddr = _T_104[4:0];
  assign mems_9_io_waddr = wptr_io_out_1[4:0];
  assign mems_9_clock = clock;
  assign mems_10_io_raddr = _T_104[4:0];
  assign mems_10_io_waddr = wptr_io_out_1[4:0];
  assign mems_10_clock = clock;
  assign mems_11_io_raddr = _T_104[4:0];
  assign mems_11_io_waddr = wptr_io_out_1[4:0];
  assign mems_11_clock = clock;
  assign mems_12_io_raddr = _T_104[4:0];
  assign mems_12_io_waddr = wptr_io_out_1[4:0];
  assign mems_12_clock = clock;
  assign mems_13_io_raddr = _T_104[4:0];
  assign mems_13_io_waddr = wptr_io_out_1[4:0];
  assign mems_13_clock = clock;
  assign mems_14_io_raddr = _T_104[4:0];
  assign mems_14_io_waddr = wptr_io_out_1[4:0];
  assign mems_14_clock = clock;
  assign mems_15_io_raddr = _T_104[4:0];
  assign mems_15_io_waddr = wptr_io_out_1[4:0];
  assign mems_15_clock = clock;
  assign FF_io_in = _T_110[3:0];
  assign FF_clock = clock;
  assign FF_reset = reset;
endmodule
module WidthConverterFIFO(
  input   clock,
  input   reset,
  input   io_enqVld,
  output  io_full,
  output  io_empty,
  output  io_almostFull
);
  wire  FIFOCore_clock;
  wire  FIFOCore_reset;
  wire  FIFOCore_io_full;
  wire  FIFOCore_io_empty;
  wire  FIFOCore_io_almostFull;
  FIFOCore_2 FIFOCore (
    .clock(FIFOCore_clock),
    .reset(FIFOCore_reset),
    .io_full(FIFOCore_io_full),
    .io_empty(FIFOCore_io_empty),
    .io_almostFull(FIFOCore_io_almostFull)
  );
  assign io_full = FIFOCore_io_full;
  assign io_empty = FIFOCore_io_empty;
  assign io_almostFull = FIFOCore_io_almostFull;
  assign FIFOCore_clock = clock;
  assign FIFOCore_reset = reset;
endmodule
module FIFOArbiterWidthConvert(
  input   clock,
  input   reset,
  output  io_empty,
  input   io_forceTag_valid,
  input   io_forceTag_bits
);
  wire  tagFF_clock;
  wire  tagFF_reset;
  wire  tagFF_io_in;
  wire  tagFF_io_out;
  wire  tagFF_io_enable;
  wire  tag;
  wire  WidthConverterFIFO_clock;
  wire  WidthConverterFIFO_reset;
  wire  WidthConverterFIFO_io_enqVld;
  wire  WidthConverterFIFO_io_full;
  wire  WidthConverterFIFO_io_empty;
  wire  WidthConverterFIFO_io_almostFull;
  wire  _T_357;
  wire  _T_358;
  FF_9 tagFF (
    .clock(tagFF_clock),
    .reset(tagFF_reset),
    .io_in(tagFF_io_in),
    .io_out(tagFF_io_out),
    .io_enable(tagFF_io_enable)
  );
  WidthConverterFIFO WidthConverterFIFO (
    .clock(WidthConverterFIFO_clock),
    .reset(WidthConverterFIFO_reset),
    .io_enqVld(WidthConverterFIFO_io_enqVld),
    .io_full(WidthConverterFIFO_io_full),
    .io_empty(WidthConverterFIFO_io_empty),
    .io_almostFull(WidthConverterFIFO_io_almostFull)
  );
  assign tag = io_forceTag_valid ? io_forceTag_bits : tagFF_io_out;
  assign _T_357 = 1'h0 == tag;
  assign _T_358 = _T_357 ? WidthConverterFIFO_io_empty : 1'h0;
  assign io_empty = _T_358;
  assign tagFF_io_in = 1'h0;
  assign tagFF_io_enable = 1'h0;
  assign tagFF_clock = clock;
  assign tagFF_reset = reset;
  assign WidthConverterFIFO_io_enqVld = 1'h0;
  assign WidthConverterFIFO_clock = clock;
  assign WidthConverterFIFO_reset = reset;
endmodule
module FF_42(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  input  [31:0] io_init,
  output [31:0] io_out,
  input         io_enable
);
  wire [31:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [31:0] RetimeWrapper_io_in;
  wire [31:0] RetimeWrapper_io_out;
  wire [31:0] _T_9;
  wire [31:0] _GEN_0;
  wire [31:0] _GEN_1;
  RetimeWrapper_1 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? io_init : _T_9;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_9;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_9 = RetimeWrapper_io_out;
endmodule
module Counter_12(
  input         clock,
  input         reset,
  input  [31:0] io_max,
  output [31:0] io_out,
  input         io_enable,
  output        io_done
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [31:0] reg$_io_in;
  wire [31:0] reg$_io_init;
  wire [31:0] reg$_io_out;
  wire  reg$_io_enable;
  wire [32:0] count;
  wire [33:0] _T_12;
  wire [32:0] newval;
  wire [32:0] _GEN_1;
  wire  isMax;
  wire [32:0] next;
  wire  _T_14;
  FF_42 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_init(reg$_io_init),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out};
  assign _T_12 = count + 33'h1;
  assign newval = _T_12[32:0];
  assign _GEN_1 = {{1'd0}, io_max};
  assign isMax = newval >= _GEN_1;
  assign next = isMax ? 33'h0 : newval;
  assign _T_14 = io_enable & isMax;
  assign io_out = count[31:0];
  assign io_done = _T_14;
  assign reg$_io_in = next[31:0];
  assign reg$_io_init = 32'h0;
  assign reg$_io_enable = io_enable;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module RetimeWrapper_43(
  input         clock,
  input         reset,
  input  [10:0] io_in,
  output [10:0] io_out
);
  wire [10:0] sr_out;
  wire [10:0] sr_in;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(11), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_44(
  input         clock,
  input         reset,
  output [10:0] io_out
);
  wire [10:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [10:0] RetimeWrapper_io_in;
  wire [10:0] RetimeWrapper_io_out;
  wire [10:0] _T_9;
  wire [10:0] _GEN_0;
  RetimeWrapper_43 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? 11'h0 : _T_9;
  assign io_out = _T_9;
  assign d = _GEN_0;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_9 = RetimeWrapper_io_out;
endmodule
module Counter_13(
  input         clock,
  input         reset,
  output [10:0] io_out
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [10:0] reg$_io_out;
  wire [11:0] count;
  FF_44 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_out(reg$_io_out)
  );
  assign count = {1'h0,reg$_io_out};
  assign io_out = count[10:0];
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module RetimeWrapper_44(
  input        clock,
  input        reset,
  input  [4:0] io_in,
  output [4:0] io_out
);
  wire [4:0] sr_out;
  wire [4:0] sr_in;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(5), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_45(
  input        clock,
  input        reset,
  input  [4:0] io_in,
  output [4:0] io_out,
  input        io_enable
);
  wire [4:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [4:0] RetimeWrapper_io_in;
  wire [4:0] RetimeWrapper_io_out;
  wire [4:0] _T_9;
  wire [4:0] _GEN_0;
  wire [4:0] _GEN_1;
  RetimeWrapper_44 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? 5'h0 : _T_9;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_9;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_9 = RetimeWrapper_io_out;
endmodule
module Counter_14(
  input   clock,
  input   reset,
  input   io_reset
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [4:0] reg$_io_in;
  wire [4:0] reg$_io_out;
  wire  reg$_io_enable;
  wire [5:0] count;
  wire [6:0] _T_12;
  wire [5:0] newval;
  wire  isMax;
  wire [5:0] next;
  wire [5:0] _GEN_0;
  FF_45 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out};
  assign _T_12 = count + 6'h1;
  assign newval = _T_12[5:0];
  assign isMax = newval >= 6'h10;
  assign next = isMax ? 6'h0 : newval;
  assign _GEN_0 = io_reset ? 6'h0 : next;
  assign reg$_io_in = _GEN_0[4:0];
  assign reg$_io_enable = io_reset;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module RetimeWrapper_557(
  input         clock,
  input         reset,
  input  [25:0] io_in,
  output [25:0] io_out
);
  wire [25:0] sr_out;
  wire [25:0] sr_in;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(26), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_558(
  input   clock,
  input   reset
);
  wire [25:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [25:0] RetimeWrapper_io_in;
  wire [25:0] RetimeWrapper_io_out;
  wire [25:0] _T_9;
  wire [25:0] _GEN_0;
  RetimeWrapper_557 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? 26'h0 : _T_9;
  assign d = _GEN_0;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_9 = RetimeWrapper_io_out;
endmodule
module SRAMByteEnable(
  input        clock,
  input  [7:0] io_wdata_0,
  input  [7:0] io_wdata_1,
  input  [7:0] io_wdata_2,
  input  [7:0] io_wdata_3,
  input  [7:0] io_wdata_4,
  input  [7:0] io_wdata_5,
  input  [7:0] io_wdata_6,
  input  [7:0] io_wdata_7,
  input  [7:0] io_wdata_8,
  input  [7:0] io_wdata_9,
  input  [7:0] io_wdata_10,
  input  [7:0] io_wdata_11,
  input  [7:0] io_wdata_12,
  input  [7:0] io_wdata_13,
  input  [7:0] io_wdata_14,
  input  [7:0] io_wdata_15,
  output [7:0] io_rdata_0,
  output [7:0] io_rdata_1,
  output [7:0] io_rdata_2,
  output [7:0] io_rdata_3,
  output [7:0] io_rdata_4,
  output [7:0] io_rdata_5,
  output [7:0] io_rdata_6,
  output [7:0] io_rdata_7,
  output [7:0] io_rdata_8,
  output [7:0] io_rdata_9,
  output [7:0] io_rdata_10,
  output [7:0] io_rdata_11,
  output [7:0] io_rdata_12,
  output [7:0] io_rdata_13,
  output [7:0] io_rdata_14,
  output [7:0] io_rdata_15
);
  reg [7:0] mem_0 [0:511];
  reg [31:0] _RAND_0;
  wire [7:0] mem_0__T_163_data;
  wire [8:0] mem_0__T_163_addr;
  wire [7:0] mem_0__T_127_data;
  wire [8:0] mem_0__T_127_addr;
  wire  mem_0__T_127_mask;
  wire  mem_0__T_127_en;
  wire  _GEN_67;
  reg [8:0] mem_0__T_163_addr_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] mem_1 [0:511];
  reg [31:0] _RAND_2;
  wire [7:0] mem_1__T_163_data;
  wire [8:0] mem_1__T_163_addr;
  wire [7:0] mem_1__T_127_data;
  wire [8:0] mem_1__T_127_addr;
  wire  mem_1__T_127_mask;
  wire  mem_1__T_127_en;
  reg [8:0] mem_1__T_163_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [7:0] mem_2 [0:511];
  reg [31:0] _RAND_4;
  wire [7:0] mem_2__T_163_data;
  wire [8:0] mem_2__T_163_addr;
  wire [7:0] mem_2__T_127_data;
  wire [8:0] mem_2__T_127_addr;
  wire  mem_2__T_127_mask;
  wire  mem_2__T_127_en;
  reg [8:0] mem_2__T_163_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [7:0] mem_3 [0:511];
  reg [31:0] _RAND_6;
  wire [7:0] mem_3__T_163_data;
  wire [8:0] mem_3__T_163_addr;
  wire [7:0] mem_3__T_127_data;
  wire [8:0] mem_3__T_127_addr;
  wire  mem_3__T_127_mask;
  wire  mem_3__T_127_en;
  reg [8:0] mem_3__T_163_addr_pipe_0;
  reg [31:0] _RAND_7;
  reg [7:0] mem_4 [0:511];
  reg [31:0] _RAND_8;
  wire [7:0] mem_4__T_163_data;
  wire [8:0] mem_4__T_163_addr;
  wire [7:0] mem_4__T_127_data;
  wire [8:0] mem_4__T_127_addr;
  wire  mem_4__T_127_mask;
  wire  mem_4__T_127_en;
  reg [8:0] mem_4__T_163_addr_pipe_0;
  reg [31:0] _RAND_9;
  reg [7:0] mem_5 [0:511];
  reg [31:0] _RAND_10;
  wire [7:0] mem_5__T_163_data;
  wire [8:0] mem_5__T_163_addr;
  wire [7:0] mem_5__T_127_data;
  wire [8:0] mem_5__T_127_addr;
  wire  mem_5__T_127_mask;
  wire  mem_5__T_127_en;
  reg [8:0] mem_5__T_163_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [7:0] mem_6 [0:511];
  reg [31:0] _RAND_12;
  wire [7:0] mem_6__T_163_data;
  wire [8:0] mem_6__T_163_addr;
  wire [7:0] mem_6__T_127_data;
  wire [8:0] mem_6__T_127_addr;
  wire  mem_6__T_127_mask;
  wire  mem_6__T_127_en;
  reg [8:0] mem_6__T_163_addr_pipe_0;
  reg [31:0] _RAND_13;
  reg [7:0] mem_7 [0:511];
  reg [31:0] _RAND_14;
  wire [7:0] mem_7__T_163_data;
  wire [8:0] mem_7__T_163_addr;
  wire [7:0] mem_7__T_127_data;
  wire [8:0] mem_7__T_127_addr;
  wire  mem_7__T_127_mask;
  wire  mem_7__T_127_en;
  reg [8:0] mem_7__T_163_addr_pipe_0;
  reg [31:0] _RAND_15;
  reg [7:0] mem_8 [0:511];
  reg [31:0] _RAND_16;
  wire [7:0] mem_8__T_163_data;
  wire [8:0] mem_8__T_163_addr;
  wire [7:0] mem_8__T_127_data;
  wire [8:0] mem_8__T_127_addr;
  wire  mem_8__T_127_mask;
  wire  mem_8__T_127_en;
  reg [8:0] mem_8__T_163_addr_pipe_0;
  reg [31:0] _RAND_17;
  reg [7:0] mem_9 [0:511];
  reg [31:0] _RAND_18;
  wire [7:0] mem_9__T_163_data;
  wire [8:0] mem_9__T_163_addr;
  wire [7:0] mem_9__T_127_data;
  wire [8:0] mem_9__T_127_addr;
  wire  mem_9__T_127_mask;
  wire  mem_9__T_127_en;
  reg [8:0] mem_9__T_163_addr_pipe_0;
  reg [31:0] _RAND_19;
  reg [7:0] mem_10 [0:511];
  reg [31:0] _RAND_20;
  wire [7:0] mem_10__T_163_data;
  wire [8:0] mem_10__T_163_addr;
  wire [7:0] mem_10__T_127_data;
  wire [8:0] mem_10__T_127_addr;
  wire  mem_10__T_127_mask;
  wire  mem_10__T_127_en;
  reg [8:0] mem_10__T_163_addr_pipe_0;
  reg [31:0] _RAND_21;
  reg [7:0] mem_11 [0:511];
  reg [31:0] _RAND_22;
  wire [7:0] mem_11__T_163_data;
  wire [8:0] mem_11__T_163_addr;
  wire [7:0] mem_11__T_127_data;
  wire [8:0] mem_11__T_127_addr;
  wire  mem_11__T_127_mask;
  wire  mem_11__T_127_en;
  reg [8:0] mem_11__T_163_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [7:0] mem_12 [0:511];
  reg [31:0] _RAND_24;
  wire [7:0] mem_12__T_163_data;
  wire [8:0] mem_12__T_163_addr;
  wire [7:0] mem_12__T_127_data;
  wire [8:0] mem_12__T_127_addr;
  wire  mem_12__T_127_mask;
  wire  mem_12__T_127_en;
  reg [8:0] mem_12__T_163_addr_pipe_0;
  reg [31:0] _RAND_25;
  reg [7:0] mem_13 [0:511];
  reg [31:0] _RAND_26;
  wire [7:0] mem_13__T_163_data;
  wire [8:0] mem_13__T_163_addr;
  wire [7:0] mem_13__T_127_data;
  wire [8:0] mem_13__T_127_addr;
  wire  mem_13__T_127_mask;
  wire  mem_13__T_127_en;
  reg [8:0] mem_13__T_163_addr_pipe_0;
  reg [31:0] _RAND_27;
  reg [7:0] mem_14 [0:511];
  reg [31:0] _RAND_28;
  wire [7:0] mem_14__T_163_data;
  wire [8:0] mem_14__T_163_addr;
  wire [7:0] mem_14__T_127_data;
  wire [8:0] mem_14__T_127_addr;
  wire  mem_14__T_127_mask;
  wire  mem_14__T_127_en;
  reg [8:0] mem_14__T_163_addr_pipe_0;
  reg [31:0] _RAND_29;
  reg [7:0] mem_15 [0:511];
  reg [31:0] _RAND_30;
  wire [7:0] mem_15__T_163_data;
  wire [8:0] mem_15__T_163_addr;
  wire [7:0] mem_15__T_127_data;
  wire [8:0] mem_15__T_127_addr;
  wire  mem_15__T_127_mask;
  wire  mem_15__T_127_en;
  reg [8:0] mem_15__T_163_addr_pipe_0;
  reg [31:0] _RAND_31;
  assign mem_0__T_163_addr = mem_0__T_163_addr_pipe_0;
  assign mem_0__T_163_data = mem_0[mem_0__T_163_addr];
  assign mem_0__T_127_data = io_wdata_0;
  assign mem_0__T_127_addr = 9'h1ff;
  assign mem_0__T_127_mask = 1'h0;
  assign mem_0__T_127_en = 1'h0;
  assign _GEN_67 = 1'h1;
  assign mem_1__T_163_addr = mem_1__T_163_addr_pipe_0;
  assign mem_1__T_163_data = mem_1[mem_1__T_163_addr];
  assign mem_1__T_127_data = io_wdata_1;
  assign mem_1__T_127_addr = 9'h1ff;
  assign mem_1__T_127_mask = 1'h0;
  assign mem_1__T_127_en = 1'h0;
  assign mem_2__T_163_addr = mem_2__T_163_addr_pipe_0;
  assign mem_2__T_163_data = mem_2[mem_2__T_163_addr];
  assign mem_2__T_127_data = io_wdata_2;
  assign mem_2__T_127_addr = 9'h1ff;
  assign mem_2__T_127_mask = 1'h0;
  assign mem_2__T_127_en = 1'h0;
  assign mem_3__T_163_addr = mem_3__T_163_addr_pipe_0;
  assign mem_3__T_163_data = mem_3[mem_3__T_163_addr];
  assign mem_3__T_127_data = io_wdata_3;
  assign mem_3__T_127_addr = 9'h1ff;
  assign mem_3__T_127_mask = 1'h0;
  assign mem_3__T_127_en = 1'h0;
  assign mem_4__T_163_addr = mem_4__T_163_addr_pipe_0;
  assign mem_4__T_163_data = mem_4[mem_4__T_163_addr];
  assign mem_4__T_127_data = io_wdata_4;
  assign mem_4__T_127_addr = 9'h1ff;
  assign mem_4__T_127_mask = 1'h0;
  assign mem_4__T_127_en = 1'h0;
  assign mem_5__T_163_addr = mem_5__T_163_addr_pipe_0;
  assign mem_5__T_163_data = mem_5[mem_5__T_163_addr];
  assign mem_5__T_127_data = io_wdata_5;
  assign mem_5__T_127_addr = 9'h1ff;
  assign mem_5__T_127_mask = 1'h0;
  assign mem_5__T_127_en = 1'h0;
  assign mem_6__T_163_addr = mem_6__T_163_addr_pipe_0;
  assign mem_6__T_163_data = mem_6[mem_6__T_163_addr];
  assign mem_6__T_127_data = io_wdata_6;
  assign mem_6__T_127_addr = 9'h1ff;
  assign mem_6__T_127_mask = 1'h0;
  assign mem_6__T_127_en = 1'h0;
  assign mem_7__T_163_addr = mem_7__T_163_addr_pipe_0;
  assign mem_7__T_163_data = mem_7[mem_7__T_163_addr];
  assign mem_7__T_127_data = io_wdata_7;
  assign mem_7__T_127_addr = 9'h1ff;
  assign mem_7__T_127_mask = 1'h0;
  assign mem_7__T_127_en = 1'h0;
  assign mem_8__T_163_addr = mem_8__T_163_addr_pipe_0;
  assign mem_8__T_163_data = mem_8[mem_8__T_163_addr];
  assign mem_8__T_127_data = io_wdata_8;
  assign mem_8__T_127_addr = 9'h1ff;
  assign mem_8__T_127_mask = 1'h0;
  assign mem_8__T_127_en = 1'h0;
  assign mem_9__T_163_addr = mem_9__T_163_addr_pipe_0;
  assign mem_9__T_163_data = mem_9[mem_9__T_163_addr];
  assign mem_9__T_127_data = io_wdata_9;
  assign mem_9__T_127_addr = 9'h1ff;
  assign mem_9__T_127_mask = 1'h0;
  assign mem_9__T_127_en = 1'h0;
  assign mem_10__T_163_addr = mem_10__T_163_addr_pipe_0;
  assign mem_10__T_163_data = mem_10[mem_10__T_163_addr];
  assign mem_10__T_127_data = io_wdata_10;
  assign mem_10__T_127_addr = 9'h1ff;
  assign mem_10__T_127_mask = 1'h0;
  assign mem_10__T_127_en = 1'h0;
  assign mem_11__T_163_addr = mem_11__T_163_addr_pipe_0;
  assign mem_11__T_163_data = mem_11[mem_11__T_163_addr];
  assign mem_11__T_127_data = io_wdata_11;
  assign mem_11__T_127_addr = 9'h1ff;
  assign mem_11__T_127_mask = 1'h0;
  assign mem_11__T_127_en = 1'h0;
  assign mem_12__T_163_addr = mem_12__T_163_addr_pipe_0;
  assign mem_12__T_163_data = mem_12[mem_12__T_163_addr];
  assign mem_12__T_127_data = io_wdata_12;
  assign mem_12__T_127_addr = 9'h1ff;
  assign mem_12__T_127_mask = 1'h0;
  assign mem_12__T_127_en = 1'h0;
  assign mem_13__T_163_addr = mem_13__T_163_addr_pipe_0;
  assign mem_13__T_163_data = mem_13[mem_13__T_163_addr];
  assign mem_13__T_127_data = io_wdata_13;
  assign mem_13__T_127_addr = 9'h1ff;
  assign mem_13__T_127_mask = 1'h0;
  assign mem_13__T_127_en = 1'h0;
  assign mem_14__T_163_addr = mem_14__T_163_addr_pipe_0;
  assign mem_14__T_163_data = mem_14[mem_14__T_163_addr];
  assign mem_14__T_127_data = io_wdata_14;
  assign mem_14__T_127_addr = 9'h1ff;
  assign mem_14__T_127_mask = 1'h0;
  assign mem_14__T_127_en = 1'h0;
  assign mem_15__T_163_addr = mem_15__T_163_addr_pipe_0;
  assign mem_15__T_163_data = mem_15[mem_15__T_163_addr];
  assign mem_15__T_127_data = io_wdata_15;
  assign mem_15__T_127_addr = 9'h1ff;
  assign mem_15__T_127_mask = 1'h0;
  assign mem_15__T_127_en = 1'h0;
  assign io_rdata_0 = mem_0__T_163_data;
  assign io_rdata_1 = mem_1__T_163_data;
  assign io_rdata_2 = mem_2__T_163_data;
  assign io_rdata_3 = mem_3__T_163_data;
  assign io_rdata_4 = mem_4__T_163_data;
  assign io_rdata_5 = mem_5__T_163_data;
  assign io_rdata_6 = mem_6__T_163_data;
  assign io_rdata_7 = mem_7__T_163_data;
  assign io_rdata_8 = mem_8__T_163_data;
  assign io_rdata_9 = mem_9__T_163_data;
  assign io_rdata_10 = mem_10__T_163_data;
  assign io_rdata_11 = mem_11__T_163_data;
  assign io_rdata_12 = mem_12__T_163_data;
  assign io_rdata_13 = mem_13__T_163_data;
  assign io_rdata_14 = mem_14__T_163_data;
  assign io_rdata_15 = mem_15__T_163_data;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_0[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem_0__T_163_addr_pipe_0 = _RAND_1[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_1[initvar] = _RAND_2[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  mem_1__T_163_addr_pipe_0 = _RAND_3[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_2[initvar] = _RAND_4[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  mem_2__T_163_addr_pipe_0 = _RAND_5[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_3[initvar] = _RAND_6[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  mem_3__T_163_addr_pipe_0 = _RAND_7[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_4[initvar] = _RAND_8[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  mem_4__T_163_addr_pipe_0 = _RAND_9[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_5[initvar] = _RAND_10[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  mem_5__T_163_addr_pipe_0 = _RAND_11[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_6[initvar] = _RAND_12[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  mem_6__T_163_addr_pipe_0 = _RAND_13[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_7[initvar] = _RAND_14[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  mem_7__T_163_addr_pipe_0 = _RAND_15[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_8[initvar] = _RAND_16[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  mem_8__T_163_addr_pipe_0 = _RAND_17[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_9[initvar] = _RAND_18[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  mem_9__T_163_addr_pipe_0 = _RAND_19[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_10[initvar] = _RAND_20[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  mem_10__T_163_addr_pipe_0 = _RAND_21[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_11[initvar] = _RAND_22[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  mem_11__T_163_addr_pipe_0 = _RAND_23[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_12[initvar] = _RAND_24[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  mem_12__T_163_addr_pipe_0 = _RAND_25[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_13[initvar] = _RAND_26[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  mem_13__T_163_addr_pipe_0 = _RAND_27[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_14[initvar] = _RAND_28[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  mem_14__T_163_addr_pipe_0 = _RAND_29[8:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    mem_15[initvar] = _RAND_30[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  mem_15__T_163_addr_pipe_0 = _RAND_31[8:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem_0__T_127_en & mem_0__T_127_mask) begin
      mem_0[mem_0__T_127_addr] <= mem_0__T_127_data;
    end
    if (_GEN_67) begin
      mem_0__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_1__T_127_en & mem_1__T_127_mask) begin
      mem_1[mem_1__T_127_addr] <= mem_1__T_127_data;
    end
    if (_GEN_67) begin
      mem_1__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_2__T_127_en & mem_2__T_127_mask) begin
      mem_2[mem_2__T_127_addr] <= mem_2__T_127_data;
    end
    if (_GEN_67) begin
      mem_2__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_3__T_127_en & mem_3__T_127_mask) begin
      mem_3[mem_3__T_127_addr] <= mem_3__T_127_data;
    end
    if (_GEN_67) begin
      mem_3__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_4__T_127_en & mem_4__T_127_mask) begin
      mem_4[mem_4__T_127_addr] <= mem_4__T_127_data;
    end
    if (_GEN_67) begin
      mem_4__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_5__T_127_en & mem_5__T_127_mask) begin
      mem_5[mem_5__T_127_addr] <= mem_5__T_127_data;
    end
    if (_GEN_67) begin
      mem_5__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_6__T_127_en & mem_6__T_127_mask) begin
      mem_6[mem_6__T_127_addr] <= mem_6__T_127_data;
    end
    if (_GEN_67) begin
      mem_6__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_7__T_127_en & mem_7__T_127_mask) begin
      mem_7[mem_7__T_127_addr] <= mem_7__T_127_data;
    end
    if (_GEN_67) begin
      mem_7__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_8__T_127_en & mem_8__T_127_mask) begin
      mem_8[mem_8__T_127_addr] <= mem_8__T_127_data;
    end
    if (_GEN_67) begin
      mem_8__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_9__T_127_en & mem_9__T_127_mask) begin
      mem_9[mem_9__T_127_addr] <= mem_9__T_127_data;
    end
    if (_GEN_67) begin
      mem_9__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_10__T_127_en & mem_10__T_127_mask) begin
      mem_10[mem_10__T_127_addr] <= mem_10__T_127_data;
    end
    if (_GEN_67) begin
      mem_10__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_11__T_127_en & mem_11__T_127_mask) begin
      mem_11[mem_11__T_127_addr] <= mem_11__T_127_data;
    end
    if (_GEN_67) begin
      mem_11__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_12__T_127_en & mem_12__T_127_mask) begin
      mem_12[mem_12__T_127_addr] <= mem_12__T_127_data;
    end
    if (_GEN_67) begin
      mem_12__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_13__T_127_en & mem_13__T_127_mask) begin
      mem_13[mem_13__T_127_addr] <= mem_13__T_127_data;
    end
    if (_GEN_67) begin
      mem_13__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_14__T_127_en & mem_14__T_127_mask) begin
      mem_14[mem_14__T_127_addr] <= mem_14__T_127_data;
    end
    if (_GEN_67) begin
      mem_14__T_163_addr_pipe_0 <= 9'h1ff;
    end
    if(mem_15__T_127_en & mem_15__T_127_mask) begin
      mem_15[mem_15__T_127_addr] <= mem_15__T_127_data;
    end
    if (_GEN_67) begin
      mem_15__T_163_addr_pipe_0 <= 9'h1ff;
    end
  end
endmodule
module CoalescingCache(
  input         clock,
  input         reset,
  output [7:0]  io_rmetaData_0,
  output [7:0]  io_rmetaData_1,
  output [7:0]  io_rmetaData_2,
  output [7:0]  io_rmetaData_3,
  output [7:0]  io_rmetaData_4,
  output [7:0]  io_rmetaData_5,
  output [7:0]  io_rmetaData_6,
  output [7:0]  io_rmetaData_7,
  output [7:0]  io_rmetaData_8,
  output [7:0]  io_rmetaData_9,
  output [7:0]  io_rmetaData_10,
  output [7:0]  io_rmetaData_11,
  output [7:0]  io_rmetaData_12,
  output [7:0]  io_rmetaData_13,
  output [7:0]  io_rmetaData_14,
  output [7:0]  io_rmetaData_15,
  input  [31:0] io_waddr,
  input  [3:0]  io_position
);
  wire  valid_0_clock;
  wire  valid_0_reset;
  wire  valid_0_io_in;
  wire  valid_0_io_out;
  wire  valid_0_io_enable;
  wire  valid_1_clock;
  wire  valid_1_reset;
  wire  valid_1_io_in;
  wire  valid_1_io_out;
  wire  valid_1_io_enable;
  wire  valid_2_clock;
  wire  valid_2_reset;
  wire  valid_2_io_in;
  wire  valid_2_io_out;
  wire  valid_2_io_enable;
  wire  valid_3_clock;
  wire  valid_3_reset;
  wire  valid_3_io_in;
  wire  valid_3_io_out;
  wire  valid_3_io_enable;
  wire  valid_4_clock;
  wire  valid_4_reset;
  wire  valid_4_io_in;
  wire  valid_4_io_out;
  wire  valid_4_io_enable;
  wire  valid_5_clock;
  wire  valid_5_reset;
  wire  valid_5_io_in;
  wire  valid_5_io_out;
  wire  valid_5_io_enable;
  wire  valid_6_clock;
  wire  valid_6_reset;
  wire  valid_6_io_in;
  wire  valid_6_io_out;
  wire  valid_6_io_enable;
  wire  valid_7_clock;
  wire  valid_7_reset;
  wire  valid_7_io_in;
  wire  valid_7_io_out;
  wire  valid_7_io_enable;
  wire  valid_8_clock;
  wire  valid_8_reset;
  wire  valid_8_io_in;
  wire  valid_8_io_out;
  wire  valid_8_io_enable;
  wire  valid_9_clock;
  wire  valid_9_reset;
  wire  valid_9_io_in;
  wire  valid_9_io_out;
  wire  valid_9_io_enable;
  wire  valid_10_clock;
  wire  valid_10_reset;
  wire  valid_10_io_in;
  wire  valid_10_io_out;
  wire  valid_10_io_enable;
  wire  valid_11_clock;
  wire  valid_11_reset;
  wire  valid_11_io_in;
  wire  valid_11_io_out;
  wire  valid_11_io_enable;
  wire  valid_12_clock;
  wire  valid_12_reset;
  wire  valid_12_io_in;
  wire  valid_12_io_out;
  wire  valid_12_io_enable;
  wire  valid_13_clock;
  wire  valid_13_reset;
  wire  valid_13_io_in;
  wire  valid_13_io_out;
  wire  valid_13_io_enable;
  wire  valid_14_clock;
  wire  valid_14_reset;
  wire  valid_14_io_in;
  wire  valid_14_io_out;
  wire  valid_14_io_enable;
  wire  valid_15_clock;
  wire  valid_15_reset;
  wire  valid_15_io_in;
  wire  valid_15_io_out;
  wire  valid_15_io_enable;
  wire  valid_16_clock;
  wire  valid_16_reset;
  wire  valid_16_io_in;
  wire  valid_16_io_out;
  wire  valid_16_io_enable;
  wire  valid_17_clock;
  wire  valid_17_reset;
  wire  valid_17_io_in;
  wire  valid_17_io_out;
  wire  valid_17_io_enable;
  wire  valid_18_clock;
  wire  valid_18_reset;
  wire  valid_18_io_in;
  wire  valid_18_io_out;
  wire  valid_18_io_enable;
  wire  valid_19_clock;
  wire  valid_19_reset;
  wire  valid_19_io_in;
  wire  valid_19_io_out;
  wire  valid_19_io_enable;
  wire  valid_20_clock;
  wire  valid_20_reset;
  wire  valid_20_io_in;
  wire  valid_20_io_out;
  wire  valid_20_io_enable;
  wire  valid_21_clock;
  wire  valid_21_reset;
  wire  valid_21_io_in;
  wire  valid_21_io_out;
  wire  valid_21_io_enable;
  wire  valid_22_clock;
  wire  valid_22_reset;
  wire  valid_22_io_in;
  wire  valid_22_io_out;
  wire  valid_22_io_enable;
  wire  valid_23_clock;
  wire  valid_23_reset;
  wire  valid_23_io_in;
  wire  valid_23_io_out;
  wire  valid_23_io_enable;
  wire  valid_24_clock;
  wire  valid_24_reset;
  wire  valid_24_io_in;
  wire  valid_24_io_out;
  wire  valid_24_io_enable;
  wire  valid_25_clock;
  wire  valid_25_reset;
  wire  valid_25_io_in;
  wire  valid_25_io_out;
  wire  valid_25_io_enable;
  wire  valid_26_clock;
  wire  valid_26_reset;
  wire  valid_26_io_in;
  wire  valid_26_io_out;
  wire  valid_26_io_enable;
  wire  valid_27_clock;
  wire  valid_27_reset;
  wire  valid_27_io_in;
  wire  valid_27_io_out;
  wire  valid_27_io_enable;
  wire  valid_28_clock;
  wire  valid_28_reset;
  wire  valid_28_io_in;
  wire  valid_28_io_out;
  wire  valid_28_io_enable;
  wire  valid_29_clock;
  wire  valid_29_reset;
  wire  valid_29_io_in;
  wire  valid_29_io_out;
  wire  valid_29_io_enable;
  wire  valid_30_clock;
  wire  valid_30_reset;
  wire  valid_30_io_in;
  wire  valid_30_io_out;
  wire  valid_30_io_enable;
  wire  valid_31_clock;
  wire  valid_31_reset;
  wire  valid_31_io_in;
  wire  valid_31_io_out;
  wire  valid_31_io_enable;
  wire  valid_32_clock;
  wire  valid_32_reset;
  wire  valid_32_io_in;
  wire  valid_32_io_out;
  wire  valid_32_io_enable;
  wire  valid_33_clock;
  wire  valid_33_reset;
  wire  valid_33_io_in;
  wire  valid_33_io_out;
  wire  valid_33_io_enable;
  wire  valid_34_clock;
  wire  valid_34_reset;
  wire  valid_34_io_in;
  wire  valid_34_io_out;
  wire  valid_34_io_enable;
  wire  valid_35_clock;
  wire  valid_35_reset;
  wire  valid_35_io_in;
  wire  valid_35_io_out;
  wire  valid_35_io_enable;
  wire  valid_36_clock;
  wire  valid_36_reset;
  wire  valid_36_io_in;
  wire  valid_36_io_out;
  wire  valid_36_io_enable;
  wire  valid_37_clock;
  wire  valid_37_reset;
  wire  valid_37_io_in;
  wire  valid_37_io_out;
  wire  valid_37_io_enable;
  wire  valid_38_clock;
  wire  valid_38_reset;
  wire  valid_38_io_in;
  wire  valid_38_io_out;
  wire  valid_38_io_enable;
  wire  valid_39_clock;
  wire  valid_39_reset;
  wire  valid_39_io_in;
  wire  valid_39_io_out;
  wire  valid_39_io_enable;
  wire  valid_40_clock;
  wire  valid_40_reset;
  wire  valid_40_io_in;
  wire  valid_40_io_out;
  wire  valid_40_io_enable;
  wire  valid_41_clock;
  wire  valid_41_reset;
  wire  valid_41_io_in;
  wire  valid_41_io_out;
  wire  valid_41_io_enable;
  wire  valid_42_clock;
  wire  valid_42_reset;
  wire  valid_42_io_in;
  wire  valid_42_io_out;
  wire  valid_42_io_enable;
  wire  valid_43_clock;
  wire  valid_43_reset;
  wire  valid_43_io_in;
  wire  valid_43_io_out;
  wire  valid_43_io_enable;
  wire  valid_44_clock;
  wire  valid_44_reset;
  wire  valid_44_io_in;
  wire  valid_44_io_out;
  wire  valid_44_io_enable;
  wire  valid_45_clock;
  wire  valid_45_reset;
  wire  valid_45_io_in;
  wire  valid_45_io_out;
  wire  valid_45_io_enable;
  wire  valid_46_clock;
  wire  valid_46_reset;
  wire  valid_46_io_in;
  wire  valid_46_io_out;
  wire  valid_46_io_enable;
  wire  valid_47_clock;
  wire  valid_47_reset;
  wire  valid_47_io_in;
  wire  valid_47_io_out;
  wire  valid_47_io_enable;
  wire  valid_48_clock;
  wire  valid_48_reset;
  wire  valid_48_io_in;
  wire  valid_48_io_out;
  wire  valid_48_io_enable;
  wire  valid_49_clock;
  wire  valid_49_reset;
  wire  valid_49_io_in;
  wire  valid_49_io_out;
  wire  valid_49_io_enable;
  wire  valid_50_clock;
  wire  valid_50_reset;
  wire  valid_50_io_in;
  wire  valid_50_io_out;
  wire  valid_50_io_enable;
  wire  valid_51_clock;
  wire  valid_51_reset;
  wire  valid_51_io_in;
  wire  valid_51_io_out;
  wire  valid_51_io_enable;
  wire  valid_52_clock;
  wire  valid_52_reset;
  wire  valid_52_io_in;
  wire  valid_52_io_out;
  wire  valid_52_io_enable;
  wire  valid_53_clock;
  wire  valid_53_reset;
  wire  valid_53_io_in;
  wire  valid_53_io_out;
  wire  valid_53_io_enable;
  wire  valid_54_clock;
  wire  valid_54_reset;
  wire  valid_54_io_in;
  wire  valid_54_io_out;
  wire  valid_54_io_enable;
  wire  valid_55_clock;
  wire  valid_55_reset;
  wire  valid_55_io_in;
  wire  valid_55_io_out;
  wire  valid_55_io_enable;
  wire  valid_56_clock;
  wire  valid_56_reset;
  wire  valid_56_io_in;
  wire  valid_56_io_out;
  wire  valid_56_io_enable;
  wire  valid_57_clock;
  wire  valid_57_reset;
  wire  valid_57_io_in;
  wire  valid_57_io_out;
  wire  valid_57_io_enable;
  wire  valid_58_clock;
  wire  valid_58_reset;
  wire  valid_58_io_in;
  wire  valid_58_io_out;
  wire  valid_58_io_enable;
  wire  valid_59_clock;
  wire  valid_59_reset;
  wire  valid_59_io_in;
  wire  valid_59_io_out;
  wire  valid_59_io_enable;
  wire  valid_60_clock;
  wire  valid_60_reset;
  wire  valid_60_io_in;
  wire  valid_60_io_out;
  wire  valid_60_io_enable;
  wire  valid_61_clock;
  wire  valid_61_reset;
  wire  valid_61_io_in;
  wire  valid_61_io_out;
  wire  valid_61_io_enable;
  wire  valid_62_clock;
  wire  valid_62_reset;
  wire  valid_62_io_in;
  wire  valid_62_io_out;
  wire  valid_62_io_enable;
  wire  valid_63_clock;
  wire  valid_63_reset;
  wire  valid_63_io_in;
  wire  valid_63_io_out;
  wire  valid_63_io_enable;
  wire  valid_64_clock;
  wire  valid_64_reset;
  wire  valid_64_io_in;
  wire  valid_64_io_out;
  wire  valid_64_io_enable;
  wire  valid_65_clock;
  wire  valid_65_reset;
  wire  valid_65_io_in;
  wire  valid_65_io_out;
  wire  valid_65_io_enable;
  wire  valid_66_clock;
  wire  valid_66_reset;
  wire  valid_66_io_in;
  wire  valid_66_io_out;
  wire  valid_66_io_enable;
  wire  valid_67_clock;
  wire  valid_67_reset;
  wire  valid_67_io_in;
  wire  valid_67_io_out;
  wire  valid_67_io_enable;
  wire  valid_68_clock;
  wire  valid_68_reset;
  wire  valid_68_io_in;
  wire  valid_68_io_out;
  wire  valid_68_io_enable;
  wire  valid_69_clock;
  wire  valid_69_reset;
  wire  valid_69_io_in;
  wire  valid_69_io_out;
  wire  valid_69_io_enable;
  wire  valid_70_clock;
  wire  valid_70_reset;
  wire  valid_70_io_in;
  wire  valid_70_io_out;
  wire  valid_70_io_enable;
  wire  valid_71_clock;
  wire  valid_71_reset;
  wire  valid_71_io_in;
  wire  valid_71_io_out;
  wire  valid_71_io_enable;
  wire  valid_72_clock;
  wire  valid_72_reset;
  wire  valid_72_io_in;
  wire  valid_72_io_out;
  wire  valid_72_io_enable;
  wire  valid_73_clock;
  wire  valid_73_reset;
  wire  valid_73_io_in;
  wire  valid_73_io_out;
  wire  valid_73_io_enable;
  wire  valid_74_clock;
  wire  valid_74_reset;
  wire  valid_74_io_in;
  wire  valid_74_io_out;
  wire  valid_74_io_enable;
  wire  valid_75_clock;
  wire  valid_75_reset;
  wire  valid_75_io_in;
  wire  valid_75_io_out;
  wire  valid_75_io_enable;
  wire  valid_76_clock;
  wire  valid_76_reset;
  wire  valid_76_io_in;
  wire  valid_76_io_out;
  wire  valid_76_io_enable;
  wire  valid_77_clock;
  wire  valid_77_reset;
  wire  valid_77_io_in;
  wire  valid_77_io_out;
  wire  valid_77_io_enable;
  wire  valid_78_clock;
  wire  valid_78_reset;
  wire  valid_78_io_in;
  wire  valid_78_io_out;
  wire  valid_78_io_enable;
  wire  valid_79_clock;
  wire  valid_79_reset;
  wire  valid_79_io_in;
  wire  valid_79_io_out;
  wire  valid_79_io_enable;
  wire  valid_80_clock;
  wire  valid_80_reset;
  wire  valid_80_io_in;
  wire  valid_80_io_out;
  wire  valid_80_io_enable;
  wire  valid_81_clock;
  wire  valid_81_reset;
  wire  valid_81_io_in;
  wire  valid_81_io_out;
  wire  valid_81_io_enable;
  wire  valid_82_clock;
  wire  valid_82_reset;
  wire  valid_82_io_in;
  wire  valid_82_io_out;
  wire  valid_82_io_enable;
  wire  valid_83_clock;
  wire  valid_83_reset;
  wire  valid_83_io_in;
  wire  valid_83_io_out;
  wire  valid_83_io_enable;
  wire  valid_84_clock;
  wire  valid_84_reset;
  wire  valid_84_io_in;
  wire  valid_84_io_out;
  wire  valid_84_io_enable;
  wire  valid_85_clock;
  wire  valid_85_reset;
  wire  valid_85_io_in;
  wire  valid_85_io_out;
  wire  valid_85_io_enable;
  wire  valid_86_clock;
  wire  valid_86_reset;
  wire  valid_86_io_in;
  wire  valid_86_io_out;
  wire  valid_86_io_enable;
  wire  valid_87_clock;
  wire  valid_87_reset;
  wire  valid_87_io_in;
  wire  valid_87_io_out;
  wire  valid_87_io_enable;
  wire  valid_88_clock;
  wire  valid_88_reset;
  wire  valid_88_io_in;
  wire  valid_88_io_out;
  wire  valid_88_io_enable;
  wire  valid_89_clock;
  wire  valid_89_reset;
  wire  valid_89_io_in;
  wire  valid_89_io_out;
  wire  valid_89_io_enable;
  wire  valid_90_clock;
  wire  valid_90_reset;
  wire  valid_90_io_in;
  wire  valid_90_io_out;
  wire  valid_90_io_enable;
  wire  valid_91_clock;
  wire  valid_91_reset;
  wire  valid_91_io_in;
  wire  valid_91_io_out;
  wire  valid_91_io_enable;
  wire  valid_92_clock;
  wire  valid_92_reset;
  wire  valid_92_io_in;
  wire  valid_92_io_out;
  wire  valid_92_io_enable;
  wire  valid_93_clock;
  wire  valid_93_reset;
  wire  valid_93_io_in;
  wire  valid_93_io_out;
  wire  valid_93_io_enable;
  wire  valid_94_clock;
  wire  valid_94_reset;
  wire  valid_94_io_in;
  wire  valid_94_io_out;
  wire  valid_94_io_enable;
  wire  valid_95_clock;
  wire  valid_95_reset;
  wire  valid_95_io_in;
  wire  valid_95_io_out;
  wire  valid_95_io_enable;
  wire  valid_96_clock;
  wire  valid_96_reset;
  wire  valid_96_io_in;
  wire  valid_96_io_out;
  wire  valid_96_io_enable;
  wire  valid_97_clock;
  wire  valid_97_reset;
  wire  valid_97_io_in;
  wire  valid_97_io_out;
  wire  valid_97_io_enable;
  wire  valid_98_clock;
  wire  valid_98_reset;
  wire  valid_98_io_in;
  wire  valid_98_io_out;
  wire  valid_98_io_enable;
  wire  valid_99_clock;
  wire  valid_99_reset;
  wire  valid_99_io_in;
  wire  valid_99_io_out;
  wire  valid_99_io_enable;
  wire  valid_100_clock;
  wire  valid_100_reset;
  wire  valid_100_io_in;
  wire  valid_100_io_out;
  wire  valid_100_io_enable;
  wire  valid_101_clock;
  wire  valid_101_reset;
  wire  valid_101_io_in;
  wire  valid_101_io_out;
  wire  valid_101_io_enable;
  wire  valid_102_clock;
  wire  valid_102_reset;
  wire  valid_102_io_in;
  wire  valid_102_io_out;
  wire  valid_102_io_enable;
  wire  valid_103_clock;
  wire  valid_103_reset;
  wire  valid_103_io_in;
  wire  valid_103_io_out;
  wire  valid_103_io_enable;
  wire  valid_104_clock;
  wire  valid_104_reset;
  wire  valid_104_io_in;
  wire  valid_104_io_out;
  wire  valid_104_io_enable;
  wire  valid_105_clock;
  wire  valid_105_reset;
  wire  valid_105_io_in;
  wire  valid_105_io_out;
  wire  valid_105_io_enable;
  wire  valid_106_clock;
  wire  valid_106_reset;
  wire  valid_106_io_in;
  wire  valid_106_io_out;
  wire  valid_106_io_enable;
  wire  valid_107_clock;
  wire  valid_107_reset;
  wire  valid_107_io_in;
  wire  valid_107_io_out;
  wire  valid_107_io_enable;
  wire  valid_108_clock;
  wire  valid_108_reset;
  wire  valid_108_io_in;
  wire  valid_108_io_out;
  wire  valid_108_io_enable;
  wire  valid_109_clock;
  wire  valid_109_reset;
  wire  valid_109_io_in;
  wire  valid_109_io_out;
  wire  valid_109_io_enable;
  wire  valid_110_clock;
  wire  valid_110_reset;
  wire  valid_110_io_in;
  wire  valid_110_io_out;
  wire  valid_110_io_enable;
  wire  valid_111_clock;
  wire  valid_111_reset;
  wire  valid_111_io_in;
  wire  valid_111_io_out;
  wire  valid_111_io_enable;
  wire  valid_112_clock;
  wire  valid_112_reset;
  wire  valid_112_io_in;
  wire  valid_112_io_out;
  wire  valid_112_io_enable;
  wire  valid_113_clock;
  wire  valid_113_reset;
  wire  valid_113_io_in;
  wire  valid_113_io_out;
  wire  valid_113_io_enable;
  wire  valid_114_clock;
  wire  valid_114_reset;
  wire  valid_114_io_in;
  wire  valid_114_io_out;
  wire  valid_114_io_enable;
  wire  valid_115_clock;
  wire  valid_115_reset;
  wire  valid_115_io_in;
  wire  valid_115_io_out;
  wire  valid_115_io_enable;
  wire  valid_116_clock;
  wire  valid_116_reset;
  wire  valid_116_io_in;
  wire  valid_116_io_out;
  wire  valid_116_io_enable;
  wire  valid_117_clock;
  wire  valid_117_reset;
  wire  valid_117_io_in;
  wire  valid_117_io_out;
  wire  valid_117_io_enable;
  wire  valid_118_clock;
  wire  valid_118_reset;
  wire  valid_118_io_in;
  wire  valid_118_io_out;
  wire  valid_118_io_enable;
  wire  valid_119_clock;
  wire  valid_119_reset;
  wire  valid_119_io_in;
  wire  valid_119_io_out;
  wire  valid_119_io_enable;
  wire  valid_120_clock;
  wire  valid_120_reset;
  wire  valid_120_io_in;
  wire  valid_120_io_out;
  wire  valid_120_io_enable;
  wire  valid_121_clock;
  wire  valid_121_reset;
  wire  valid_121_io_in;
  wire  valid_121_io_out;
  wire  valid_121_io_enable;
  wire  valid_122_clock;
  wire  valid_122_reset;
  wire  valid_122_io_in;
  wire  valid_122_io_out;
  wire  valid_122_io_enable;
  wire  valid_123_clock;
  wire  valid_123_reset;
  wire  valid_123_io_in;
  wire  valid_123_io_out;
  wire  valid_123_io_enable;
  wire  valid_124_clock;
  wire  valid_124_reset;
  wire  valid_124_io_in;
  wire  valid_124_io_out;
  wire  valid_124_io_enable;
  wire  valid_125_clock;
  wire  valid_125_reset;
  wire  valid_125_io_in;
  wire  valid_125_io_out;
  wire  valid_125_io_enable;
  wire  valid_126_clock;
  wire  valid_126_reset;
  wire  valid_126_io_in;
  wire  valid_126_io_out;
  wire  valid_126_io_enable;
  wire  valid_127_clock;
  wire  valid_127_reset;
  wire  valid_127_io_in;
  wire  valid_127_io_out;
  wire  valid_127_io_enable;
  wire  valid_128_clock;
  wire  valid_128_reset;
  wire  valid_128_io_in;
  wire  valid_128_io_out;
  wire  valid_128_io_enable;
  wire  valid_129_clock;
  wire  valid_129_reset;
  wire  valid_129_io_in;
  wire  valid_129_io_out;
  wire  valid_129_io_enable;
  wire  valid_130_clock;
  wire  valid_130_reset;
  wire  valid_130_io_in;
  wire  valid_130_io_out;
  wire  valid_130_io_enable;
  wire  valid_131_clock;
  wire  valid_131_reset;
  wire  valid_131_io_in;
  wire  valid_131_io_out;
  wire  valid_131_io_enable;
  wire  valid_132_clock;
  wire  valid_132_reset;
  wire  valid_132_io_in;
  wire  valid_132_io_out;
  wire  valid_132_io_enable;
  wire  valid_133_clock;
  wire  valid_133_reset;
  wire  valid_133_io_in;
  wire  valid_133_io_out;
  wire  valid_133_io_enable;
  wire  valid_134_clock;
  wire  valid_134_reset;
  wire  valid_134_io_in;
  wire  valid_134_io_out;
  wire  valid_134_io_enable;
  wire  valid_135_clock;
  wire  valid_135_reset;
  wire  valid_135_io_in;
  wire  valid_135_io_out;
  wire  valid_135_io_enable;
  wire  valid_136_clock;
  wire  valid_136_reset;
  wire  valid_136_io_in;
  wire  valid_136_io_out;
  wire  valid_136_io_enable;
  wire  valid_137_clock;
  wire  valid_137_reset;
  wire  valid_137_io_in;
  wire  valid_137_io_out;
  wire  valid_137_io_enable;
  wire  valid_138_clock;
  wire  valid_138_reset;
  wire  valid_138_io_in;
  wire  valid_138_io_out;
  wire  valid_138_io_enable;
  wire  valid_139_clock;
  wire  valid_139_reset;
  wire  valid_139_io_in;
  wire  valid_139_io_out;
  wire  valid_139_io_enable;
  wire  valid_140_clock;
  wire  valid_140_reset;
  wire  valid_140_io_in;
  wire  valid_140_io_out;
  wire  valid_140_io_enable;
  wire  valid_141_clock;
  wire  valid_141_reset;
  wire  valid_141_io_in;
  wire  valid_141_io_out;
  wire  valid_141_io_enable;
  wire  valid_142_clock;
  wire  valid_142_reset;
  wire  valid_142_io_in;
  wire  valid_142_io_out;
  wire  valid_142_io_enable;
  wire  valid_143_clock;
  wire  valid_143_reset;
  wire  valid_143_io_in;
  wire  valid_143_io_out;
  wire  valid_143_io_enable;
  wire  valid_144_clock;
  wire  valid_144_reset;
  wire  valid_144_io_in;
  wire  valid_144_io_out;
  wire  valid_144_io_enable;
  wire  valid_145_clock;
  wire  valid_145_reset;
  wire  valid_145_io_in;
  wire  valid_145_io_out;
  wire  valid_145_io_enable;
  wire  valid_146_clock;
  wire  valid_146_reset;
  wire  valid_146_io_in;
  wire  valid_146_io_out;
  wire  valid_146_io_enable;
  wire  valid_147_clock;
  wire  valid_147_reset;
  wire  valid_147_io_in;
  wire  valid_147_io_out;
  wire  valid_147_io_enable;
  wire  valid_148_clock;
  wire  valid_148_reset;
  wire  valid_148_io_in;
  wire  valid_148_io_out;
  wire  valid_148_io_enable;
  wire  valid_149_clock;
  wire  valid_149_reset;
  wire  valid_149_io_in;
  wire  valid_149_io_out;
  wire  valid_149_io_enable;
  wire  valid_150_clock;
  wire  valid_150_reset;
  wire  valid_150_io_in;
  wire  valid_150_io_out;
  wire  valid_150_io_enable;
  wire  valid_151_clock;
  wire  valid_151_reset;
  wire  valid_151_io_in;
  wire  valid_151_io_out;
  wire  valid_151_io_enable;
  wire  valid_152_clock;
  wire  valid_152_reset;
  wire  valid_152_io_in;
  wire  valid_152_io_out;
  wire  valid_152_io_enable;
  wire  valid_153_clock;
  wire  valid_153_reset;
  wire  valid_153_io_in;
  wire  valid_153_io_out;
  wire  valid_153_io_enable;
  wire  valid_154_clock;
  wire  valid_154_reset;
  wire  valid_154_io_in;
  wire  valid_154_io_out;
  wire  valid_154_io_enable;
  wire  valid_155_clock;
  wire  valid_155_reset;
  wire  valid_155_io_in;
  wire  valid_155_io_out;
  wire  valid_155_io_enable;
  wire  valid_156_clock;
  wire  valid_156_reset;
  wire  valid_156_io_in;
  wire  valid_156_io_out;
  wire  valid_156_io_enable;
  wire  valid_157_clock;
  wire  valid_157_reset;
  wire  valid_157_io_in;
  wire  valid_157_io_out;
  wire  valid_157_io_enable;
  wire  valid_158_clock;
  wire  valid_158_reset;
  wire  valid_158_io_in;
  wire  valid_158_io_out;
  wire  valid_158_io_enable;
  wire  valid_159_clock;
  wire  valid_159_reset;
  wire  valid_159_io_in;
  wire  valid_159_io_out;
  wire  valid_159_io_enable;
  wire  valid_160_clock;
  wire  valid_160_reset;
  wire  valid_160_io_in;
  wire  valid_160_io_out;
  wire  valid_160_io_enable;
  wire  valid_161_clock;
  wire  valid_161_reset;
  wire  valid_161_io_in;
  wire  valid_161_io_out;
  wire  valid_161_io_enable;
  wire  valid_162_clock;
  wire  valid_162_reset;
  wire  valid_162_io_in;
  wire  valid_162_io_out;
  wire  valid_162_io_enable;
  wire  valid_163_clock;
  wire  valid_163_reset;
  wire  valid_163_io_in;
  wire  valid_163_io_out;
  wire  valid_163_io_enable;
  wire  valid_164_clock;
  wire  valid_164_reset;
  wire  valid_164_io_in;
  wire  valid_164_io_out;
  wire  valid_164_io_enable;
  wire  valid_165_clock;
  wire  valid_165_reset;
  wire  valid_165_io_in;
  wire  valid_165_io_out;
  wire  valid_165_io_enable;
  wire  valid_166_clock;
  wire  valid_166_reset;
  wire  valid_166_io_in;
  wire  valid_166_io_out;
  wire  valid_166_io_enable;
  wire  valid_167_clock;
  wire  valid_167_reset;
  wire  valid_167_io_in;
  wire  valid_167_io_out;
  wire  valid_167_io_enable;
  wire  valid_168_clock;
  wire  valid_168_reset;
  wire  valid_168_io_in;
  wire  valid_168_io_out;
  wire  valid_168_io_enable;
  wire  valid_169_clock;
  wire  valid_169_reset;
  wire  valid_169_io_in;
  wire  valid_169_io_out;
  wire  valid_169_io_enable;
  wire  valid_170_clock;
  wire  valid_170_reset;
  wire  valid_170_io_in;
  wire  valid_170_io_out;
  wire  valid_170_io_enable;
  wire  valid_171_clock;
  wire  valid_171_reset;
  wire  valid_171_io_in;
  wire  valid_171_io_out;
  wire  valid_171_io_enable;
  wire  valid_172_clock;
  wire  valid_172_reset;
  wire  valid_172_io_in;
  wire  valid_172_io_out;
  wire  valid_172_io_enable;
  wire  valid_173_clock;
  wire  valid_173_reset;
  wire  valid_173_io_in;
  wire  valid_173_io_out;
  wire  valid_173_io_enable;
  wire  valid_174_clock;
  wire  valid_174_reset;
  wire  valid_174_io_in;
  wire  valid_174_io_out;
  wire  valid_174_io_enable;
  wire  valid_175_clock;
  wire  valid_175_reset;
  wire  valid_175_io_in;
  wire  valid_175_io_out;
  wire  valid_175_io_enable;
  wire  valid_176_clock;
  wire  valid_176_reset;
  wire  valid_176_io_in;
  wire  valid_176_io_out;
  wire  valid_176_io_enable;
  wire  valid_177_clock;
  wire  valid_177_reset;
  wire  valid_177_io_in;
  wire  valid_177_io_out;
  wire  valid_177_io_enable;
  wire  valid_178_clock;
  wire  valid_178_reset;
  wire  valid_178_io_in;
  wire  valid_178_io_out;
  wire  valid_178_io_enable;
  wire  valid_179_clock;
  wire  valid_179_reset;
  wire  valid_179_io_in;
  wire  valid_179_io_out;
  wire  valid_179_io_enable;
  wire  valid_180_clock;
  wire  valid_180_reset;
  wire  valid_180_io_in;
  wire  valid_180_io_out;
  wire  valid_180_io_enable;
  wire  valid_181_clock;
  wire  valid_181_reset;
  wire  valid_181_io_in;
  wire  valid_181_io_out;
  wire  valid_181_io_enable;
  wire  valid_182_clock;
  wire  valid_182_reset;
  wire  valid_182_io_in;
  wire  valid_182_io_out;
  wire  valid_182_io_enable;
  wire  valid_183_clock;
  wire  valid_183_reset;
  wire  valid_183_io_in;
  wire  valid_183_io_out;
  wire  valid_183_io_enable;
  wire  valid_184_clock;
  wire  valid_184_reset;
  wire  valid_184_io_in;
  wire  valid_184_io_out;
  wire  valid_184_io_enable;
  wire  valid_185_clock;
  wire  valid_185_reset;
  wire  valid_185_io_in;
  wire  valid_185_io_out;
  wire  valid_185_io_enable;
  wire  valid_186_clock;
  wire  valid_186_reset;
  wire  valid_186_io_in;
  wire  valid_186_io_out;
  wire  valid_186_io_enable;
  wire  valid_187_clock;
  wire  valid_187_reset;
  wire  valid_187_io_in;
  wire  valid_187_io_out;
  wire  valid_187_io_enable;
  wire  valid_188_clock;
  wire  valid_188_reset;
  wire  valid_188_io_in;
  wire  valid_188_io_out;
  wire  valid_188_io_enable;
  wire  valid_189_clock;
  wire  valid_189_reset;
  wire  valid_189_io_in;
  wire  valid_189_io_out;
  wire  valid_189_io_enable;
  wire  valid_190_clock;
  wire  valid_190_reset;
  wire  valid_190_io_in;
  wire  valid_190_io_out;
  wire  valid_190_io_enable;
  wire  valid_191_clock;
  wire  valid_191_reset;
  wire  valid_191_io_in;
  wire  valid_191_io_out;
  wire  valid_191_io_enable;
  wire  valid_192_clock;
  wire  valid_192_reset;
  wire  valid_192_io_in;
  wire  valid_192_io_out;
  wire  valid_192_io_enable;
  wire  valid_193_clock;
  wire  valid_193_reset;
  wire  valid_193_io_in;
  wire  valid_193_io_out;
  wire  valid_193_io_enable;
  wire  valid_194_clock;
  wire  valid_194_reset;
  wire  valid_194_io_in;
  wire  valid_194_io_out;
  wire  valid_194_io_enable;
  wire  valid_195_clock;
  wire  valid_195_reset;
  wire  valid_195_io_in;
  wire  valid_195_io_out;
  wire  valid_195_io_enable;
  wire  valid_196_clock;
  wire  valid_196_reset;
  wire  valid_196_io_in;
  wire  valid_196_io_out;
  wire  valid_196_io_enable;
  wire  valid_197_clock;
  wire  valid_197_reset;
  wire  valid_197_io_in;
  wire  valid_197_io_out;
  wire  valid_197_io_enable;
  wire  valid_198_clock;
  wire  valid_198_reset;
  wire  valid_198_io_in;
  wire  valid_198_io_out;
  wire  valid_198_io_enable;
  wire  valid_199_clock;
  wire  valid_199_reset;
  wire  valid_199_io_in;
  wire  valid_199_io_out;
  wire  valid_199_io_enable;
  wire  valid_200_clock;
  wire  valid_200_reset;
  wire  valid_200_io_in;
  wire  valid_200_io_out;
  wire  valid_200_io_enable;
  wire  valid_201_clock;
  wire  valid_201_reset;
  wire  valid_201_io_in;
  wire  valid_201_io_out;
  wire  valid_201_io_enable;
  wire  valid_202_clock;
  wire  valid_202_reset;
  wire  valid_202_io_in;
  wire  valid_202_io_out;
  wire  valid_202_io_enable;
  wire  valid_203_clock;
  wire  valid_203_reset;
  wire  valid_203_io_in;
  wire  valid_203_io_out;
  wire  valid_203_io_enable;
  wire  valid_204_clock;
  wire  valid_204_reset;
  wire  valid_204_io_in;
  wire  valid_204_io_out;
  wire  valid_204_io_enable;
  wire  valid_205_clock;
  wire  valid_205_reset;
  wire  valid_205_io_in;
  wire  valid_205_io_out;
  wire  valid_205_io_enable;
  wire  valid_206_clock;
  wire  valid_206_reset;
  wire  valid_206_io_in;
  wire  valid_206_io_out;
  wire  valid_206_io_enable;
  wire  valid_207_clock;
  wire  valid_207_reset;
  wire  valid_207_io_in;
  wire  valid_207_io_out;
  wire  valid_207_io_enable;
  wire  valid_208_clock;
  wire  valid_208_reset;
  wire  valid_208_io_in;
  wire  valid_208_io_out;
  wire  valid_208_io_enable;
  wire  valid_209_clock;
  wire  valid_209_reset;
  wire  valid_209_io_in;
  wire  valid_209_io_out;
  wire  valid_209_io_enable;
  wire  valid_210_clock;
  wire  valid_210_reset;
  wire  valid_210_io_in;
  wire  valid_210_io_out;
  wire  valid_210_io_enable;
  wire  valid_211_clock;
  wire  valid_211_reset;
  wire  valid_211_io_in;
  wire  valid_211_io_out;
  wire  valid_211_io_enable;
  wire  valid_212_clock;
  wire  valid_212_reset;
  wire  valid_212_io_in;
  wire  valid_212_io_out;
  wire  valid_212_io_enable;
  wire  valid_213_clock;
  wire  valid_213_reset;
  wire  valid_213_io_in;
  wire  valid_213_io_out;
  wire  valid_213_io_enable;
  wire  valid_214_clock;
  wire  valid_214_reset;
  wire  valid_214_io_in;
  wire  valid_214_io_out;
  wire  valid_214_io_enable;
  wire  valid_215_clock;
  wire  valid_215_reset;
  wire  valid_215_io_in;
  wire  valid_215_io_out;
  wire  valid_215_io_enable;
  wire  valid_216_clock;
  wire  valid_216_reset;
  wire  valid_216_io_in;
  wire  valid_216_io_out;
  wire  valid_216_io_enable;
  wire  valid_217_clock;
  wire  valid_217_reset;
  wire  valid_217_io_in;
  wire  valid_217_io_out;
  wire  valid_217_io_enable;
  wire  valid_218_clock;
  wire  valid_218_reset;
  wire  valid_218_io_in;
  wire  valid_218_io_out;
  wire  valid_218_io_enable;
  wire  valid_219_clock;
  wire  valid_219_reset;
  wire  valid_219_io_in;
  wire  valid_219_io_out;
  wire  valid_219_io_enable;
  wire  valid_220_clock;
  wire  valid_220_reset;
  wire  valid_220_io_in;
  wire  valid_220_io_out;
  wire  valid_220_io_enable;
  wire  valid_221_clock;
  wire  valid_221_reset;
  wire  valid_221_io_in;
  wire  valid_221_io_out;
  wire  valid_221_io_enable;
  wire  valid_222_clock;
  wire  valid_222_reset;
  wire  valid_222_io_in;
  wire  valid_222_io_out;
  wire  valid_222_io_enable;
  wire  valid_223_clock;
  wire  valid_223_reset;
  wire  valid_223_io_in;
  wire  valid_223_io_out;
  wire  valid_223_io_enable;
  wire  valid_224_clock;
  wire  valid_224_reset;
  wire  valid_224_io_in;
  wire  valid_224_io_out;
  wire  valid_224_io_enable;
  wire  valid_225_clock;
  wire  valid_225_reset;
  wire  valid_225_io_in;
  wire  valid_225_io_out;
  wire  valid_225_io_enable;
  wire  valid_226_clock;
  wire  valid_226_reset;
  wire  valid_226_io_in;
  wire  valid_226_io_out;
  wire  valid_226_io_enable;
  wire  valid_227_clock;
  wire  valid_227_reset;
  wire  valid_227_io_in;
  wire  valid_227_io_out;
  wire  valid_227_io_enable;
  wire  valid_228_clock;
  wire  valid_228_reset;
  wire  valid_228_io_in;
  wire  valid_228_io_out;
  wire  valid_228_io_enable;
  wire  valid_229_clock;
  wire  valid_229_reset;
  wire  valid_229_io_in;
  wire  valid_229_io_out;
  wire  valid_229_io_enable;
  wire  valid_230_clock;
  wire  valid_230_reset;
  wire  valid_230_io_in;
  wire  valid_230_io_out;
  wire  valid_230_io_enable;
  wire  valid_231_clock;
  wire  valid_231_reset;
  wire  valid_231_io_in;
  wire  valid_231_io_out;
  wire  valid_231_io_enable;
  wire  valid_232_clock;
  wire  valid_232_reset;
  wire  valid_232_io_in;
  wire  valid_232_io_out;
  wire  valid_232_io_enable;
  wire  valid_233_clock;
  wire  valid_233_reset;
  wire  valid_233_io_in;
  wire  valid_233_io_out;
  wire  valid_233_io_enable;
  wire  valid_234_clock;
  wire  valid_234_reset;
  wire  valid_234_io_in;
  wire  valid_234_io_out;
  wire  valid_234_io_enable;
  wire  valid_235_clock;
  wire  valid_235_reset;
  wire  valid_235_io_in;
  wire  valid_235_io_out;
  wire  valid_235_io_enable;
  wire  valid_236_clock;
  wire  valid_236_reset;
  wire  valid_236_io_in;
  wire  valid_236_io_out;
  wire  valid_236_io_enable;
  wire  valid_237_clock;
  wire  valid_237_reset;
  wire  valid_237_io_in;
  wire  valid_237_io_out;
  wire  valid_237_io_enable;
  wire  valid_238_clock;
  wire  valid_238_reset;
  wire  valid_238_io_in;
  wire  valid_238_io_out;
  wire  valid_238_io_enable;
  wire  valid_239_clock;
  wire  valid_239_reset;
  wire  valid_239_io_in;
  wire  valid_239_io_out;
  wire  valid_239_io_enable;
  wire  valid_240_clock;
  wire  valid_240_reset;
  wire  valid_240_io_in;
  wire  valid_240_io_out;
  wire  valid_240_io_enable;
  wire  valid_241_clock;
  wire  valid_241_reset;
  wire  valid_241_io_in;
  wire  valid_241_io_out;
  wire  valid_241_io_enable;
  wire  valid_242_clock;
  wire  valid_242_reset;
  wire  valid_242_io_in;
  wire  valid_242_io_out;
  wire  valid_242_io_enable;
  wire  valid_243_clock;
  wire  valid_243_reset;
  wire  valid_243_io_in;
  wire  valid_243_io_out;
  wire  valid_243_io_enable;
  wire  valid_244_clock;
  wire  valid_244_reset;
  wire  valid_244_io_in;
  wire  valid_244_io_out;
  wire  valid_244_io_enable;
  wire  valid_245_clock;
  wire  valid_245_reset;
  wire  valid_245_io_in;
  wire  valid_245_io_out;
  wire  valid_245_io_enable;
  wire  valid_246_clock;
  wire  valid_246_reset;
  wire  valid_246_io_in;
  wire  valid_246_io_out;
  wire  valid_246_io_enable;
  wire  valid_247_clock;
  wire  valid_247_reset;
  wire  valid_247_io_in;
  wire  valid_247_io_out;
  wire  valid_247_io_enable;
  wire  valid_248_clock;
  wire  valid_248_reset;
  wire  valid_248_io_in;
  wire  valid_248_io_out;
  wire  valid_248_io_enable;
  wire  valid_249_clock;
  wire  valid_249_reset;
  wire  valid_249_io_in;
  wire  valid_249_io_out;
  wire  valid_249_io_enable;
  wire  valid_250_clock;
  wire  valid_250_reset;
  wire  valid_250_io_in;
  wire  valid_250_io_out;
  wire  valid_250_io_enable;
  wire  valid_251_clock;
  wire  valid_251_reset;
  wire  valid_251_io_in;
  wire  valid_251_io_out;
  wire  valid_251_io_enable;
  wire  valid_252_clock;
  wire  valid_252_reset;
  wire  valid_252_io_in;
  wire  valid_252_io_out;
  wire  valid_252_io_enable;
  wire  valid_253_clock;
  wire  valid_253_reset;
  wire  valid_253_io_in;
  wire  valid_253_io_out;
  wire  valid_253_io_enable;
  wire  valid_254_clock;
  wire  valid_254_reset;
  wire  valid_254_io_in;
  wire  valid_254_io_out;
  wire  valid_254_io_enable;
  wire  valid_255_clock;
  wire  valid_255_reset;
  wire  valid_255_io_in;
  wire  valid_255_io_out;
  wire  valid_255_io_enable;
  wire  valid_256_clock;
  wire  valid_256_reset;
  wire  valid_256_io_in;
  wire  valid_256_io_out;
  wire  valid_256_io_enable;
  wire  valid_257_clock;
  wire  valid_257_reset;
  wire  valid_257_io_in;
  wire  valid_257_io_out;
  wire  valid_257_io_enable;
  wire  valid_258_clock;
  wire  valid_258_reset;
  wire  valid_258_io_in;
  wire  valid_258_io_out;
  wire  valid_258_io_enable;
  wire  valid_259_clock;
  wire  valid_259_reset;
  wire  valid_259_io_in;
  wire  valid_259_io_out;
  wire  valid_259_io_enable;
  wire  valid_260_clock;
  wire  valid_260_reset;
  wire  valid_260_io_in;
  wire  valid_260_io_out;
  wire  valid_260_io_enable;
  wire  valid_261_clock;
  wire  valid_261_reset;
  wire  valid_261_io_in;
  wire  valid_261_io_out;
  wire  valid_261_io_enable;
  wire  valid_262_clock;
  wire  valid_262_reset;
  wire  valid_262_io_in;
  wire  valid_262_io_out;
  wire  valid_262_io_enable;
  wire  valid_263_clock;
  wire  valid_263_reset;
  wire  valid_263_io_in;
  wire  valid_263_io_out;
  wire  valid_263_io_enable;
  wire  valid_264_clock;
  wire  valid_264_reset;
  wire  valid_264_io_in;
  wire  valid_264_io_out;
  wire  valid_264_io_enable;
  wire  valid_265_clock;
  wire  valid_265_reset;
  wire  valid_265_io_in;
  wire  valid_265_io_out;
  wire  valid_265_io_enable;
  wire  valid_266_clock;
  wire  valid_266_reset;
  wire  valid_266_io_in;
  wire  valid_266_io_out;
  wire  valid_266_io_enable;
  wire  valid_267_clock;
  wire  valid_267_reset;
  wire  valid_267_io_in;
  wire  valid_267_io_out;
  wire  valid_267_io_enable;
  wire  valid_268_clock;
  wire  valid_268_reset;
  wire  valid_268_io_in;
  wire  valid_268_io_out;
  wire  valid_268_io_enable;
  wire  valid_269_clock;
  wire  valid_269_reset;
  wire  valid_269_io_in;
  wire  valid_269_io_out;
  wire  valid_269_io_enable;
  wire  valid_270_clock;
  wire  valid_270_reset;
  wire  valid_270_io_in;
  wire  valid_270_io_out;
  wire  valid_270_io_enable;
  wire  valid_271_clock;
  wire  valid_271_reset;
  wire  valid_271_io_in;
  wire  valid_271_io_out;
  wire  valid_271_io_enable;
  wire  valid_272_clock;
  wire  valid_272_reset;
  wire  valid_272_io_in;
  wire  valid_272_io_out;
  wire  valid_272_io_enable;
  wire  valid_273_clock;
  wire  valid_273_reset;
  wire  valid_273_io_in;
  wire  valid_273_io_out;
  wire  valid_273_io_enable;
  wire  valid_274_clock;
  wire  valid_274_reset;
  wire  valid_274_io_in;
  wire  valid_274_io_out;
  wire  valid_274_io_enable;
  wire  valid_275_clock;
  wire  valid_275_reset;
  wire  valid_275_io_in;
  wire  valid_275_io_out;
  wire  valid_275_io_enable;
  wire  valid_276_clock;
  wire  valid_276_reset;
  wire  valid_276_io_in;
  wire  valid_276_io_out;
  wire  valid_276_io_enable;
  wire  valid_277_clock;
  wire  valid_277_reset;
  wire  valid_277_io_in;
  wire  valid_277_io_out;
  wire  valid_277_io_enable;
  wire  valid_278_clock;
  wire  valid_278_reset;
  wire  valid_278_io_in;
  wire  valid_278_io_out;
  wire  valid_278_io_enable;
  wire  valid_279_clock;
  wire  valid_279_reset;
  wire  valid_279_io_in;
  wire  valid_279_io_out;
  wire  valid_279_io_enable;
  wire  valid_280_clock;
  wire  valid_280_reset;
  wire  valid_280_io_in;
  wire  valid_280_io_out;
  wire  valid_280_io_enable;
  wire  valid_281_clock;
  wire  valid_281_reset;
  wire  valid_281_io_in;
  wire  valid_281_io_out;
  wire  valid_281_io_enable;
  wire  valid_282_clock;
  wire  valid_282_reset;
  wire  valid_282_io_in;
  wire  valid_282_io_out;
  wire  valid_282_io_enable;
  wire  valid_283_clock;
  wire  valid_283_reset;
  wire  valid_283_io_in;
  wire  valid_283_io_out;
  wire  valid_283_io_enable;
  wire  valid_284_clock;
  wire  valid_284_reset;
  wire  valid_284_io_in;
  wire  valid_284_io_out;
  wire  valid_284_io_enable;
  wire  valid_285_clock;
  wire  valid_285_reset;
  wire  valid_285_io_in;
  wire  valid_285_io_out;
  wire  valid_285_io_enable;
  wire  valid_286_clock;
  wire  valid_286_reset;
  wire  valid_286_io_in;
  wire  valid_286_io_out;
  wire  valid_286_io_enable;
  wire  valid_287_clock;
  wire  valid_287_reset;
  wire  valid_287_io_in;
  wire  valid_287_io_out;
  wire  valid_287_io_enable;
  wire  valid_288_clock;
  wire  valid_288_reset;
  wire  valid_288_io_in;
  wire  valid_288_io_out;
  wire  valid_288_io_enable;
  wire  valid_289_clock;
  wire  valid_289_reset;
  wire  valid_289_io_in;
  wire  valid_289_io_out;
  wire  valid_289_io_enable;
  wire  valid_290_clock;
  wire  valid_290_reset;
  wire  valid_290_io_in;
  wire  valid_290_io_out;
  wire  valid_290_io_enable;
  wire  valid_291_clock;
  wire  valid_291_reset;
  wire  valid_291_io_in;
  wire  valid_291_io_out;
  wire  valid_291_io_enable;
  wire  valid_292_clock;
  wire  valid_292_reset;
  wire  valid_292_io_in;
  wire  valid_292_io_out;
  wire  valid_292_io_enable;
  wire  valid_293_clock;
  wire  valid_293_reset;
  wire  valid_293_io_in;
  wire  valid_293_io_out;
  wire  valid_293_io_enable;
  wire  valid_294_clock;
  wire  valid_294_reset;
  wire  valid_294_io_in;
  wire  valid_294_io_out;
  wire  valid_294_io_enable;
  wire  valid_295_clock;
  wire  valid_295_reset;
  wire  valid_295_io_in;
  wire  valid_295_io_out;
  wire  valid_295_io_enable;
  wire  valid_296_clock;
  wire  valid_296_reset;
  wire  valid_296_io_in;
  wire  valid_296_io_out;
  wire  valid_296_io_enable;
  wire  valid_297_clock;
  wire  valid_297_reset;
  wire  valid_297_io_in;
  wire  valid_297_io_out;
  wire  valid_297_io_enable;
  wire  valid_298_clock;
  wire  valid_298_reset;
  wire  valid_298_io_in;
  wire  valid_298_io_out;
  wire  valid_298_io_enable;
  wire  valid_299_clock;
  wire  valid_299_reset;
  wire  valid_299_io_in;
  wire  valid_299_io_out;
  wire  valid_299_io_enable;
  wire  valid_300_clock;
  wire  valid_300_reset;
  wire  valid_300_io_in;
  wire  valid_300_io_out;
  wire  valid_300_io_enable;
  wire  valid_301_clock;
  wire  valid_301_reset;
  wire  valid_301_io_in;
  wire  valid_301_io_out;
  wire  valid_301_io_enable;
  wire  valid_302_clock;
  wire  valid_302_reset;
  wire  valid_302_io_in;
  wire  valid_302_io_out;
  wire  valid_302_io_enable;
  wire  valid_303_clock;
  wire  valid_303_reset;
  wire  valid_303_io_in;
  wire  valid_303_io_out;
  wire  valid_303_io_enable;
  wire  valid_304_clock;
  wire  valid_304_reset;
  wire  valid_304_io_in;
  wire  valid_304_io_out;
  wire  valid_304_io_enable;
  wire  valid_305_clock;
  wire  valid_305_reset;
  wire  valid_305_io_in;
  wire  valid_305_io_out;
  wire  valid_305_io_enable;
  wire  valid_306_clock;
  wire  valid_306_reset;
  wire  valid_306_io_in;
  wire  valid_306_io_out;
  wire  valid_306_io_enable;
  wire  valid_307_clock;
  wire  valid_307_reset;
  wire  valid_307_io_in;
  wire  valid_307_io_out;
  wire  valid_307_io_enable;
  wire  valid_308_clock;
  wire  valid_308_reset;
  wire  valid_308_io_in;
  wire  valid_308_io_out;
  wire  valid_308_io_enable;
  wire  valid_309_clock;
  wire  valid_309_reset;
  wire  valid_309_io_in;
  wire  valid_309_io_out;
  wire  valid_309_io_enable;
  wire  valid_310_clock;
  wire  valid_310_reset;
  wire  valid_310_io_in;
  wire  valid_310_io_out;
  wire  valid_310_io_enable;
  wire  valid_311_clock;
  wire  valid_311_reset;
  wire  valid_311_io_in;
  wire  valid_311_io_out;
  wire  valid_311_io_enable;
  wire  valid_312_clock;
  wire  valid_312_reset;
  wire  valid_312_io_in;
  wire  valid_312_io_out;
  wire  valid_312_io_enable;
  wire  valid_313_clock;
  wire  valid_313_reset;
  wire  valid_313_io_in;
  wire  valid_313_io_out;
  wire  valid_313_io_enable;
  wire  valid_314_clock;
  wire  valid_314_reset;
  wire  valid_314_io_in;
  wire  valid_314_io_out;
  wire  valid_314_io_enable;
  wire  valid_315_clock;
  wire  valid_315_reset;
  wire  valid_315_io_in;
  wire  valid_315_io_out;
  wire  valid_315_io_enable;
  wire  valid_316_clock;
  wire  valid_316_reset;
  wire  valid_316_io_in;
  wire  valid_316_io_out;
  wire  valid_316_io_enable;
  wire  valid_317_clock;
  wire  valid_317_reset;
  wire  valid_317_io_in;
  wire  valid_317_io_out;
  wire  valid_317_io_enable;
  wire  valid_318_clock;
  wire  valid_318_reset;
  wire  valid_318_io_in;
  wire  valid_318_io_out;
  wire  valid_318_io_enable;
  wire  valid_319_clock;
  wire  valid_319_reset;
  wire  valid_319_io_in;
  wire  valid_319_io_out;
  wire  valid_319_io_enable;
  wire  valid_320_clock;
  wire  valid_320_reset;
  wire  valid_320_io_in;
  wire  valid_320_io_out;
  wire  valid_320_io_enable;
  wire  valid_321_clock;
  wire  valid_321_reset;
  wire  valid_321_io_in;
  wire  valid_321_io_out;
  wire  valid_321_io_enable;
  wire  valid_322_clock;
  wire  valid_322_reset;
  wire  valid_322_io_in;
  wire  valid_322_io_out;
  wire  valid_322_io_enable;
  wire  valid_323_clock;
  wire  valid_323_reset;
  wire  valid_323_io_in;
  wire  valid_323_io_out;
  wire  valid_323_io_enable;
  wire  valid_324_clock;
  wire  valid_324_reset;
  wire  valid_324_io_in;
  wire  valid_324_io_out;
  wire  valid_324_io_enable;
  wire  valid_325_clock;
  wire  valid_325_reset;
  wire  valid_325_io_in;
  wire  valid_325_io_out;
  wire  valid_325_io_enable;
  wire  valid_326_clock;
  wire  valid_326_reset;
  wire  valid_326_io_in;
  wire  valid_326_io_out;
  wire  valid_326_io_enable;
  wire  valid_327_clock;
  wire  valid_327_reset;
  wire  valid_327_io_in;
  wire  valid_327_io_out;
  wire  valid_327_io_enable;
  wire  valid_328_clock;
  wire  valid_328_reset;
  wire  valid_328_io_in;
  wire  valid_328_io_out;
  wire  valid_328_io_enable;
  wire  valid_329_clock;
  wire  valid_329_reset;
  wire  valid_329_io_in;
  wire  valid_329_io_out;
  wire  valid_329_io_enable;
  wire  valid_330_clock;
  wire  valid_330_reset;
  wire  valid_330_io_in;
  wire  valid_330_io_out;
  wire  valid_330_io_enable;
  wire  valid_331_clock;
  wire  valid_331_reset;
  wire  valid_331_io_in;
  wire  valid_331_io_out;
  wire  valid_331_io_enable;
  wire  valid_332_clock;
  wire  valid_332_reset;
  wire  valid_332_io_in;
  wire  valid_332_io_out;
  wire  valid_332_io_enable;
  wire  valid_333_clock;
  wire  valid_333_reset;
  wire  valid_333_io_in;
  wire  valid_333_io_out;
  wire  valid_333_io_enable;
  wire  valid_334_clock;
  wire  valid_334_reset;
  wire  valid_334_io_in;
  wire  valid_334_io_out;
  wire  valid_334_io_enable;
  wire  valid_335_clock;
  wire  valid_335_reset;
  wire  valid_335_io_in;
  wire  valid_335_io_out;
  wire  valid_335_io_enable;
  wire  valid_336_clock;
  wire  valid_336_reset;
  wire  valid_336_io_in;
  wire  valid_336_io_out;
  wire  valid_336_io_enable;
  wire  valid_337_clock;
  wire  valid_337_reset;
  wire  valid_337_io_in;
  wire  valid_337_io_out;
  wire  valid_337_io_enable;
  wire  valid_338_clock;
  wire  valid_338_reset;
  wire  valid_338_io_in;
  wire  valid_338_io_out;
  wire  valid_338_io_enable;
  wire  valid_339_clock;
  wire  valid_339_reset;
  wire  valid_339_io_in;
  wire  valid_339_io_out;
  wire  valid_339_io_enable;
  wire  valid_340_clock;
  wire  valid_340_reset;
  wire  valid_340_io_in;
  wire  valid_340_io_out;
  wire  valid_340_io_enable;
  wire  valid_341_clock;
  wire  valid_341_reset;
  wire  valid_341_io_in;
  wire  valid_341_io_out;
  wire  valid_341_io_enable;
  wire  valid_342_clock;
  wire  valid_342_reset;
  wire  valid_342_io_in;
  wire  valid_342_io_out;
  wire  valid_342_io_enable;
  wire  valid_343_clock;
  wire  valid_343_reset;
  wire  valid_343_io_in;
  wire  valid_343_io_out;
  wire  valid_343_io_enable;
  wire  valid_344_clock;
  wire  valid_344_reset;
  wire  valid_344_io_in;
  wire  valid_344_io_out;
  wire  valid_344_io_enable;
  wire  valid_345_clock;
  wire  valid_345_reset;
  wire  valid_345_io_in;
  wire  valid_345_io_out;
  wire  valid_345_io_enable;
  wire  valid_346_clock;
  wire  valid_346_reset;
  wire  valid_346_io_in;
  wire  valid_346_io_out;
  wire  valid_346_io_enable;
  wire  valid_347_clock;
  wire  valid_347_reset;
  wire  valid_347_io_in;
  wire  valid_347_io_out;
  wire  valid_347_io_enable;
  wire  valid_348_clock;
  wire  valid_348_reset;
  wire  valid_348_io_in;
  wire  valid_348_io_out;
  wire  valid_348_io_enable;
  wire  valid_349_clock;
  wire  valid_349_reset;
  wire  valid_349_io_in;
  wire  valid_349_io_out;
  wire  valid_349_io_enable;
  wire  valid_350_clock;
  wire  valid_350_reset;
  wire  valid_350_io_in;
  wire  valid_350_io_out;
  wire  valid_350_io_enable;
  wire  valid_351_clock;
  wire  valid_351_reset;
  wire  valid_351_io_in;
  wire  valid_351_io_out;
  wire  valid_351_io_enable;
  wire  valid_352_clock;
  wire  valid_352_reset;
  wire  valid_352_io_in;
  wire  valid_352_io_out;
  wire  valid_352_io_enable;
  wire  valid_353_clock;
  wire  valid_353_reset;
  wire  valid_353_io_in;
  wire  valid_353_io_out;
  wire  valid_353_io_enable;
  wire  valid_354_clock;
  wire  valid_354_reset;
  wire  valid_354_io_in;
  wire  valid_354_io_out;
  wire  valid_354_io_enable;
  wire  valid_355_clock;
  wire  valid_355_reset;
  wire  valid_355_io_in;
  wire  valid_355_io_out;
  wire  valid_355_io_enable;
  wire  valid_356_clock;
  wire  valid_356_reset;
  wire  valid_356_io_in;
  wire  valid_356_io_out;
  wire  valid_356_io_enable;
  wire  valid_357_clock;
  wire  valid_357_reset;
  wire  valid_357_io_in;
  wire  valid_357_io_out;
  wire  valid_357_io_enable;
  wire  valid_358_clock;
  wire  valid_358_reset;
  wire  valid_358_io_in;
  wire  valid_358_io_out;
  wire  valid_358_io_enable;
  wire  valid_359_clock;
  wire  valid_359_reset;
  wire  valid_359_io_in;
  wire  valid_359_io_out;
  wire  valid_359_io_enable;
  wire  valid_360_clock;
  wire  valid_360_reset;
  wire  valid_360_io_in;
  wire  valid_360_io_out;
  wire  valid_360_io_enable;
  wire  valid_361_clock;
  wire  valid_361_reset;
  wire  valid_361_io_in;
  wire  valid_361_io_out;
  wire  valid_361_io_enable;
  wire  valid_362_clock;
  wire  valid_362_reset;
  wire  valid_362_io_in;
  wire  valid_362_io_out;
  wire  valid_362_io_enable;
  wire  valid_363_clock;
  wire  valid_363_reset;
  wire  valid_363_io_in;
  wire  valid_363_io_out;
  wire  valid_363_io_enable;
  wire  valid_364_clock;
  wire  valid_364_reset;
  wire  valid_364_io_in;
  wire  valid_364_io_out;
  wire  valid_364_io_enable;
  wire  valid_365_clock;
  wire  valid_365_reset;
  wire  valid_365_io_in;
  wire  valid_365_io_out;
  wire  valid_365_io_enable;
  wire  valid_366_clock;
  wire  valid_366_reset;
  wire  valid_366_io_in;
  wire  valid_366_io_out;
  wire  valid_366_io_enable;
  wire  valid_367_clock;
  wire  valid_367_reset;
  wire  valid_367_io_in;
  wire  valid_367_io_out;
  wire  valid_367_io_enable;
  wire  valid_368_clock;
  wire  valid_368_reset;
  wire  valid_368_io_in;
  wire  valid_368_io_out;
  wire  valid_368_io_enable;
  wire  valid_369_clock;
  wire  valid_369_reset;
  wire  valid_369_io_in;
  wire  valid_369_io_out;
  wire  valid_369_io_enable;
  wire  valid_370_clock;
  wire  valid_370_reset;
  wire  valid_370_io_in;
  wire  valid_370_io_out;
  wire  valid_370_io_enable;
  wire  valid_371_clock;
  wire  valid_371_reset;
  wire  valid_371_io_in;
  wire  valid_371_io_out;
  wire  valid_371_io_enable;
  wire  valid_372_clock;
  wire  valid_372_reset;
  wire  valid_372_io_in;
  wire  valid_372_io_out;
  wire  valid_372_io_enable;
  wire  valid_373_clock;
  wire  valid_373_reset;
  wire  valid_373_io_in;
  wire  valid_373_io_out;
  wire  valid_373_io_enable;
  wire  valid_374_clock;
  wire  valid_374_reset;
  wire  valid_374_io_in;
  wire  valid_374_io_out;
  wire  valid_374_io_enable;
  wire  valid_375_clock;
  wire  valid_375_reset;
  wire  valid_375_io_in;
  wire  valid_375_io_out;
  wire  valid_375_io_enable;
  wire  valid_376_clock;
  wire  valid_376_reset;
  wire  valid_376_io_in;
  wire  valid_376_io_out;
  wire  valid_376_io_enable;
  wire  valid_377_clock;
  wire  valid_377_reset;
  wire  valid_377_io_in;
  wire  valid_377_io_out;
  wire  valid_377_io_enable;
  wire  valid_378_clock;
  wire  valid_378_reset;
  wire  valid_378_io_in;
  wire  valid_378_io_out;
  wire  valid_378_io_enable;
  wire  valid_379_clock;
  wire  valid_379_reset;
  wire  valid_379_io_in;
  wire  valid_379_io_out;
  wire  valid_379_io_enable;
  wire  valid_380_clock;
  wire  valid_380_reset;
  wire  valid_380_io_in;
  wire  valid_380_io_out;
  wire  valid_380_io_enable;
  wire  valid_381_clock;
  wire  valid_381_reset;
  wire  valid_381_io_in;
  wire  valid_381_io_out;
  wire  valid_381_io_enable;
  wire  valid_382_clock;
  wire  valid_382_reset;
  wire  valid_382_io_in;
  wire  valid_382_io_out;
  wire  valid_382_io_enable;
  wire  valid_383_clock;
  wire  valid_383_reset;
  wire  valid_383_io_in;
  wire  valid_383_io_out;
  wire  valid_383_io_enable;
  wire  valid_384_clock;
  wire  valid_384_reset;
  wire  valid_384_io_in;
  wire  valid_384_io_out;
  wire  valid_384_io_enable;
  wire  valid_385_clock;
  wire  valid_385_reset;
  wire  valid_385_io_in;
  wire  valid_385_io_out;
  wire  valid_385_io_enable;
  wire  valid_386_clock;
  wire  valid_386_reset;
  wire  valid_386_io_in;
  wire  valid_386_io_out;
  wire  valid_386_io_enable;
  wire  valid_387_clock;
  wire  valid_387_reset;
  wire  valid_387_io_in;
  wire  valid_387_io_out;
  wire  valid_387_io_enable;
  wire  valid_388_clock;
  wire  valid_388_reset;
  wire  valid_388_io_in;
  wire  valid_388_io_out;
  wire  valid_388_io_enable;
  wire  valid_389_clock;
  wire  valid_389_reset;
  wire  valid_389_io_in;
  wire  valid_389_io_out;
  wire  valid_389_io_enable;
  wire  valid_390_clock;
  wire  valid_390_reset;
  wire  valid_390_io_in;
  wire  valid_390_io_out;
  wire  valid_390_io_enable;
  wire  valid_391_clock;
  wire  valid_391_reset;
  wire  valid_391_io_in;
  wire  valid_391_io_out;
  wire  valid_391_io_enable;
  wire  valid_392_clock;
  wire  valid_392_reset;
  wire  valid_392_io_in;
  wire  valid_392_io_out;
  wire  valid_392_io_enable;
  wire  valid_393_clock;
  wire  valid_393_reset;
  wire  valid_393_io_in;
  wire  valid_393_io_out;
  wire  valid_393_io_enable;
  wire  valid_394_clock;
  wire  valid_394_reset;
  wire  valid_394_io_in;
  wire  valid_394_io_out;
  wire  valid_394_io_enable;
  wire  valid_395_clock;
  wire  valid_395_reset;
  wire  valid_395_io_in;
  wire  valid_395_io_out;
  wire  valid_395_io_enable;
  wire  valid_396_clock;
  wire  valid_396_reset;
  wire  valid_396_io_in;
  wire  valid_396_io_out;
  wire  valid_396_io_enable;
  wire  valid_397_clock;
  wire  valid_397_reset;
  wire  valid_397_io_in;
  wire  valid_397_io_out;
  wire  valid_397_io_enable;
  wire  valid_398_clock;
  wire  valid_398_reset;
  wire  valid_398_io_in;
  wire  valid_398_io_out;
  wire  valid_398_io_enable;
  wire  valid_399_clock;
  wire  valid_399_reset;
  wire  valid_399_io_in;
  wire  valid_399_io_out;
  wire  valid_399_io_enable;
  wire  valid_400_clock;
  wire  valid_400_reset;
  wire  valid_400_io_in;
  wire  valid_400_io_out;
  wire  valid_400_io_enable;
  wire  valid_401_clock;
  wire  valid_401_reset;
  wire  valid_401_io_in;
  wire  valid_401_io_out;
  wire  valid_401_io_enable;
  wire  valid_402_clock;
  wire  valid_402_reset;
  wire  valid_402_io_in;
  wire  valid_402_io_out;
  wire  valid_402_io_enable;
  wire  valid_403_clock;
  wire  valid_403_reset;
  wire  valid_403_io_in;
  wire  valid_403_io_out;
  wire  valid_403_io_enable;
  wire  valid_404_clock;
  wire  valid_404_reset;
  wire  valid_404_io_in;
  wire  valid_404_io_out;
  wire  valid_404_io_enable;
  wire  valid_405_clock;
  wire  valid_405_reset;
  wire  valid_405_io_in;
  wire  valid_405_io_out;
  wire  valid_405_io_enable;
  wire  valid_406_clock;
  wire  valid_406_reset;
  wire  valid_406_io_in;
  wire  valid_406_io_out;
  wire  valid_406_io_enable;
  wire  valid_407_clock;
  wire  valid_407_reset;
  wire  valid_407_io_in;
  wire  valid_407_io_out;
  wire  valid_407_io_enable;
  wire  valid_408_clock;
  wire  valid_408_reset;
  wire  valid_408_io_in;
  wire  valid_408_io_out;
  wire  valid_408_io_enable;
  wire  valid_409_clock;
  wire  valid_409_reset;
  wire  valid_409_io_in;
  wire  valid_409_io_out;
  wire  valid_409_io_enable;
  wire  valid_410_clock;
  wire  valid_410_reset;
  wire  valid_410_io_in;
  wire  valid_410_io_out;
  wire  valid_410_io_enable;
  wire  valid_411_clock;
  wire  valid_411_reset;
  wire  valid_411_io_in;
  wire  valid_411_io_out;
  wire  valid_411_io_enable;
  wire  valid_412_clock;
  wire  valid_412_reset;
  wire  valid_412_io_in;
  wire  valid_412_io_out;
  wire  valid_412_io_enable;
  wire  valid_413_clock;
  wire  valid_413_reset;
  wire  valid_413_io_in;
  wire  valid_413_io_out;
  wire  valid_413_io_enable;
  wire  valid_414_clock;
  wire  valid_414_reset;
  wire  valid_414_io_in;
  wire  valid_414_io_out;
  wire  valid_414_io_enable;
  wire  valid_415_clock;
  wire  valid_415_reset;
  wire  valid_415_io_in;
  wire  valid_415_io_out;
  wire  valid_415_io_enable;
  wire  valid_416_clock;
  wire  valid_416_reset;
  wire  valid_416_io_in;
  wire  valid_416_io_out;
  wire  valid_416_io_enable;
  wire  valid_417_clock;
  wire  valid_417_reset;
  wire  valid_417_io_in;
  wire  valid_417_io_out;
  wire  valid_417_io_enable;
  wire  valid_418_clock;
  wire  valid_418_reset;
  wire  valid_418_io_in;
  wire  valid_418_io_out;
  wire  valid_418_io_enable;
  wire  valid_419_clock;
  wire  valid_419_reset;
  wire  valid_419_io_in;
  wire  valid_419_io_out;
  wire  valid_419_io_enable;
  wire  valid_420_clock;
  wire  valid_420_reset;
  wire  valid_420_io_in;
  wire  valid_420_io_out;
  wire  valid_420_io_enable;
  wire  valid_421_clock;
  wire  valid_421_reset;
  wire  valid_421_io_in;
  wire  valid_421_io_out;
  wire  valid_421_io_enable;
  wire  valid_422_clock;
  wire  valid_422_reset;
  wire  valid_422_io_in;
  wire  valid_422_io_out;
  wire  valid_422_io_enable;
  wire  valid_423_clock;
  wire  valid_423_reset;
  wire  valid_423_io_in;
  wire  valid_423_io_out;
  wire  valid_423_io_enable;
  wire  valid_424_clock;
  wire  valid_424_reset;
  wire  valid_424_io_in;
  wire  valid_424_io_out;
  wire  valid_424_io_enable;
  wire  valid_425_clock;
  wire  valid_425_reset;
  wire  valid_425_io_in;
  wire  valid_425_io_out;
  wire  valid_425_io_enable;
  wire  valid_426_clock;
  wire  valid_426_reset;
  wire  valid_426_io_in;
  wire  valid_426_io_out;
  wire  valid_426_io_enable;
  wire  valid_427_clock;
  wire  valid_427_reset;
  wire  valid_427_io_in;
  wire  valid_427_io_out;
  wire  valid_427_io_enable;
  wire  valid_428_clock;
  wire  valid_428_reset;
  wire  valid_428_io_in;
  wire  valid_428_io_out;
  wire  valid_428_io_enable;
  wire  valid_429_clock;
  wire  valid_429_reset;
  wire  valid_429_io_in;
  wire  valid_429_io_out;
  wire  valid_429_io_enable;
  wire  valid_430_clock;
  wire  valid_430_reset;
  wire  valid_430_io_in;
  wire  valid_430_io_out;
  wire  valid_430_io_enable;
  wire  valid_431_clock;
  wire  valid_431_reset;
  wire  valid_431_io_in;
  wire  valid_431_io_out;
  wire  valid_431_io_enable;
  wire  valid_432_clock;
  wire  valid_432_reset;
  wire  valid_432_io_in;
  wire  valid_432_io_out;
  wire  valid_432_io_enable;
  wire  valid_433_clock;
  wire  valid_433_reset;
  wire  valid_433_io_in;
  wire  valid_433_io_out;
  wire  valid_433_io_enable;
  wire  valid_434_clock;
  wire  valid_434_reset;
  wire  valid_434_io_in;
  wire  valid_434_io_out;
  wire  valid_434_io_enable;
  wire  valid_435_clock;
  wire  valid_435_reset;
  wire  valid_435_io_in;
  wire  valid_435_io_out;
  wire  valid_435_io_enable;
  wire  valid_436_clock;
  wire  valid_436_reset;
  wire  valid_436_io_in;
  wire  valid_436_io_out;
  wire  valid_436_io_enable;
  wire  valid_437_clock;
  wire  valid_437_reset;
  wire  valid_437_io_in;
  wire  valid_437_io_out;
  wire  valid_437_io_enable;
  wire  valid_438_clock;
  wire  valid_438_reset;
  wire  valid_438_io_in;
  wire  valid_438_io_out;
  wire  valid_438_io_enable;
  wire  valid_439_clock;
  wire  valid_439_reset;
  wire  valid_439_io_in;
  wire  valid_439_io_out;
  wire  valid_439_io_enable;
  wire  valid_440_clock;
  wire  valid_440_reset;
  wire  valid_440_io_in;
  wire  valid_440_io_out;
  wire  valid_440_io_enable;
  wire  valid_441_clock;
  wire  valid_441_reset;
  wire  valid_441_io_in;
  wire  valid_441_io_out;
  wire  valid_441_io_enable;
  wire  valid_442_clock;
  wire  valid_442_reset;
  wire  valid_442_io_in;
  wire  valid_442_io_out;
  wire  valid_442_io_enable;
  wire  valid_443_clock;
  wire  valid_443_reset;
  wire  valid_443_io_in;
  wire  valid_443_io_out;
  wire  valid_443_io_enable;
  wire  valid_444_clock;
  wire  valid_444_reset;
  wire  valid_444_io_in;
  wire  valid_444_io_out;
  wire  valid_444_io_enable;
  wire  valid_445_clock;
  wire  valid_445_reset;
  wire  valid_445_io_in;
  wire  valid_445_io_out;
  wire  valid_445_io_enable;
  wire  valid_446_clock;
  wire  valid_446_reset;
  wire  valid_446_io_in;
  wire  valid_446_io_out;
  wire  valid_446_io_enable;
  wire  valid_447_clock;
  wire  valid_447_reset;
  wire  valid_447_io_in;
  wire  valid_447_io_out;
  wire  valid_447_io_enable;
  wire  valid_448_clock;
  wire  valid_448_reset;
  wire  valid_448_io_in;
  wire  valid_448_io_out;
  wire  valid_448_io_enable;
  wire  valid_449_clock;
  wire  valid_449_reset;
  wire  valid_449_io_in;
  wire  valid_449_io_out;
  wire  valid_449_io_enable;
  wire  valid_450_clock;
  wire  valid_450_reset;
  wire  valid_450_io_in;
  wire  valid_450_io_out;
  wire  valid_450_io_enable;
  wire  valid_451_clock;
  wire  valid_451_reset;
  wire  valid_451_io_in;
  wire  valid_451_io_out;
  wire  valid_451_io_enable;
  wire  valid_452_clock;
  wire  valid_452_reset;
  wire  valid_452_io_in;
  wire  valid_452_io_out;
  wire  valid_452_io_enable;
  wire  valid_453_clock;
  wire  valid_453_reset;
  wire  valid_453_io_in;
  wire  valid_453_io_out;
  wire  valid_453_io_enable;
  wire  valid_454_clock;
  wire  valid_454_reset;
  wire  valid_454_io_in;
  wire  valid_454_io_out;
  wire  valid_454_io_enable;
  wire  valid_455_clock;
  wire  valid_455_reset;
  wire  valid_455_io_in;
  wire  valid_455_io_out;
  wire  valid_455_io_enable;
  wire  valid_456_clock;
  wire  valid_456_reset;
  wire  valid_456_io_in;
  wire  valid_456_io_out;
  wire  valid_456_io_enable;
  wire  valid_457_clock;
  wire  valid_457_reset;
  wire  valid_457_io_in;
  wire  valid_457_io_out;
  wire  valid_457_io_enable;
  wire  valid_458_clock;
  wire  valid_458_reset;
  wire  valid_458_io_in;
  wire  valid_458_io_out;
  wire  valid_458_io_enable;
  wire  valid_459_clock;
  wire  valid_459_reset;
  wire  valid_459_io_in;
  wire  valid_459_io_out;
  wire  valid_459_io_enable;
  wire  valid_460_clock;
  wire  valid_460_reset;
  wire  valid_460_io_in;
  wire  valid_460_io_out;
  wire  valid_460_io_enable;
  wire  valid_461_clock;
  wire  valid_461_reset;
  wire  valid_461_io_in;
  wire  valid_461_io_out;
  wire  valid_461_io_enable;
  wire  valid_462_clock;
  wire  valid_462_reset;
  wire  valid_462_io_in;
  wire  valid_462_io_out;
  wire  valid_462_io_enable;
  wire  valid_463_clock;
  wire  valid_463_reset;
  wire  valid_463_io_in;
  wire  valid_463_io_out;
  wire  valid_463_io_enable;
  wire  valid_464_clock;
  wire  valid_464_reset;
  wire  valid_464_io_in;
  wire  valid_464_io_out;
  wire  valid_464_io_enable;
  wire  valid_465_clock;
  wire  valid_465_reset;
  wire  valid_465_io_in;
  wire  valid_465_io_out;
  wire  valid_465_io_enable;
  wire  valid_466_clock;
  wire  valid_466_reset;
  wire  valid_466_io_in;
  wire  valid_466_io_out;
  wire  valid_466_io_enable;
  wire  valid_467_clock;
  wire  valid_467_reset;
  wire  valid_467_io_in;
  wire  valid_467_io_out;
  wire  valid_467_io_enable;
  wire  valid_468_clock;
  wire  valid_468_reset;
  wire  valid_468_io_in;
  wire  valid_468_io_out;
  wire  valid_468_io_enable;
  wire  valid_469_clock;
  wire  valid_469_reset;
  wire  valid_469_io_in;
  wire  valid_469_io_out;
  wire  valid_469_io_enable;
  wire  valid_470_clock;
  wire  valid_470_reset;
  wire  valid_470_io_in;
  wire  valid_470_io_out;
  wire  valid_470_io_enable;
  wire  valid_471_clock;
  wire  valid_471_reset;
  wire  valid_471_io_in;
  wire  valid_471_io_out;
  wire  valid_471_io_enable;
  wire  valid_472_clock;
  wire  valid_472_reset;
  wire  valid_472_io_in;
  wire  valid_472_io_out;
  wire  valid_472_io_enable;
  wire  valid_473_clock;
  wire  valid_473_reset;
  wire  valid_473_io_in;
  wire  valid_473_io_out;
  wire  valid_473_io_enable;
  wire  valid_474_clock;
  wire  valid_474_reset;
  wire  valid_474_io_in;
  wire  valid_474_io_out;
  wire  valid_474_io_enable;
  wire  valid_475_clock;
  wire  valid_475_reset;
  wire  valid_475_io_in;
  wire  valid_475_io_out;
  wire  valid_475_io_enable;
  wire  valid_476_clock;
  wire  valid_476_reset;
  wire  valid_476_io_in;
  wire  valid_476_io_out;
  wire  valid_476_io_enable;
  wire  valid_477_clock;
  wire  valid_477_reset;
  wire  valid_477_io_in;
  wire  valid_477_io_out;
  wire  valid_477_io_enable;
  wire  valid_478_clock;
  wire  valid_478_reset;
  wire  valid_478_io_in;
  wire  valid_478_io_out;
  wire  valid_478_io_enable;
  wire  valid_479_clock;
  wire  valid_479_reset;
  wire  valid_479_io_in;
  wire  valid_479_io_out;
  wire  valid_479_io_enable;
  wire  valid_480_clock;
  wire  valid_480_reset;
  wire  valid_480_io_in;
  wire  valid_480_io_out;
  wire  valid_480_io_enable;
  wire  valid_481_clock;
  wire  valid_481_reset;
  wire  valid_481_io_in;
  wire  valid_481_io_out;
  wire  valid_481_io_enable;
  wire  valid_482_clock;
  wire  valid_482_reset;
  wire  valid_482_io_in;
  wire  valid_482_io_out;
  wire  valid_482_io_enable;
  wire  valid_483_clock;
  wire  valid_483_reset;
  wire  valid_483_io_in;
  wire  valid_483_io_out;
  wire  valid_483_io_enable;
  wire  valid_484_clock;
  wire  valid_484_reset;
  wire  valid_484_io_in;
  wire  valid_484_io_out;
  wire  valid_484_io_enable;
  wire  valid_485_clock;
  wire  valid_485_reset;
  wire  valid_485_io_in;
  wire  valid_485_io_out;
  wire  valid_485_io_enable;
  wire  valid_486_clock;
  wire  valid_486_reset;
  wire  valid_486_io_in;
  wire  valid_486_io_out;
  wire  valid_486_io_enable;
  wire  valid_487_clock;
  wire  valid_487_reset;
  wire  valid_487_io_in;
  wire  valid_487_io_out;
  wire  valid_487_io_enable;
  wire  valid_488_clock;
  wire  valid_488_reset;
  wire  valid_488_io_in;
  wire  valid_488_io_out;
  wire  valid_488_io_enable;
  wire  valid_489_clock;
  wire  valid_489_reset;
  wire  valid_489_io_in;
  wire  valid_489_io_out;
  wire  valid_489_io_enable;
  wire  valid_490_clock;
  wire  valid_490_reset;
  wire  valid_490_io_in;
  wire  valid_490_io_out;
  wire  valid_490_io_enable;
  wire  valid_491_clock;
  wire  valid_491_reset;
  wire  valid_491_io_in;
  wire  valid_491_io_out;
  wire  valid_491_io_enable;
  wire  valid_492_clock;
  wire  valid_492_reset;
  wire  valid_492_io_in;
  wire  valid_492_io_out;
  wire  valid_492_io_enable;
  wire  valid_493_clock;
  wire  valid_493_reset;
  wire  valid_493_io_in;
  wire  valid_493_io_out;
  wire  valid_493_io_enable;
  wire  valid_494_clock;
  wire  valid_494_reset;
  wire  valid_494_io_in;
  wire  valid_494_io_out;
  wire  valid_494_io_enable;
  wire  valid_495_clock;
  wire  valid_495_reset;
  wire  valid_495_io_in;
  wire  valid_495_io_out;
  wire  valid_495_io_enable;
  wire  valid_496_clock;
  wire  valid_496_reset;
  wire  valid_496_io_in;
  wire  valid_496_io_out;
  wire  valid_496_io_enable;
  wire  valid_497_clock;
  wire  valid_497_reset;
  wire  valid_497_io_in;
  wire  valid_497_io_out;
  wire  valid_497_io_enable;
  wire  valid_498_clock;
  wire  valid_498_reset;
  wire  valid_498_io_in;
  wire  valid_498_io_out;
  wire  valid_498_io_enable;
  wire  valid_499_clock;
  wire  valid_499_reset;
  wire  valid_499_io_in;
  wire  valid_499_io_out;
  wire  valid_499_io_enable;
  wire  valid_500_clock;
  wire  valid_500_reset;
  wire  valid_500_io_in;
  wire  valid_500_io_out;
  wire  valid_500_io_enable;
  wire  valid_501_clock;
  wire  valid_501_reset;
  wire  valid_501_io_in;
  wire  valid_501_io_out;
  wire  valid_501_io_enable;
  wire  valid_502_clock;
  wire  valid_502_reset;
  wire  valid_502_io_in;
  wire  valid_502_io_out;
  wire  valid_502_io_enable;
  wire  valid_503_clock;
  wire  valid_503_reset;
  wire  valid_503_io_in;
  wire  valid_503_io_out;
  wire  valid_503_io_enable;
  wire  valid_504_clock;
  wire  valid_504_reset;
  wire  valid_504_io_in;
  wire  valid_504_io_out;
  wire  valid_504_io_enable;
  wire  valid_505_clock;
  wire  valid_505_reset;
  wire  valid_505_io_in;
  wire  valid_505_io_out;
  wire  valid_505_io_enable;
  wire  valid_506_clock;
  wire  valid_506_reset;
  wire  valid_506_io_in;
  wire  valid_506_io_out;
  wire  valid_506_io_enable;
  wire  valid_507_clock;
  wire  valid_507_reset;
  wire  valid_507_io_in;
  wire  valid_507_io_out;
  wire  valid_507_io_enable;
  wire  valid_508_clock;
  wire  valid_508_reset;
  wire  valid_508_io_in;
  wire  valid_508_io_out;
  wire  valid_508_io_enable;
  wire  valid_509_clock;
  wire  valid_509_reset;
  wire  valid_509_io_in;
  wire  valid_509_io_out;
  wire  valid_509_io_enable;
  wire  valid_510_clock;
  wire  valid_510_reset;
  wire  valid_510_io_in;
  wire  valid_510_io_out;
  wire  valid_510_io_enable;
  wire  valid_511_clock;
  wire  valid_511_reset;
  wire  valid_511_io_in;
  wire  valid_511_io_out;
  wire  valid_511_io_enable;
  wire  tags_0_clock;
  wire  tags_0_reset;
  wire  tags_1_clock;
  wire  tags_1_reset;
  wire  tags_2_clock;
  wire  tags_2_reset;
  wire  tags_3_clock;
  wire  tags_3_reset;
  wire  tags_4_clock;
  wire  tags_4_reset;
  wire  tags_5_clock;
  wire  tags_5_reset;
  wire  tags_6_clock;
  wire  tags_6_reset;
  wire  tags_7_clock;
  wire  tags_7_reset;
  wire  tags_8_clock;
  wire  tags_8_reset;
  wire  tags_9_clock;
  wire  tags_9_reset;
  wire  tags_10_clock;
  wire  tags_10_reset;
  wire  tags_11_clock;
  wire  tags_11_reset;
  wire  tags_12_clock;
  wire  tags_12_reset;
  wire  tags_13_clock;
  wire  tags_13_reset;
  wire  tags_14_clock;
  wire  tags_14_reset;
  wire  tags_15_clock;
  wire  tags_15_reset;
  wire  tags_16_clock;
  wire  tags_16_reset;
  wire  tags_17_clock;
  wire  tags_17_reset;
  wire  tags_18_clock;
  wire  tags_18_reset;
  wire  tags_19_clock;
  wire  tags_19_reset;
  wire  tags_20_clock;
  wire  tags_20_reset;
  wire  tags_21_clock;
  wire  tags_21_reset;
  wire  tags_22_clock;
  wire  tags_22_reset;
  wire  tags_23_clock;
  wire  tags_23_reset;
  wire  tags_24_clock;
  wire  tags_24_reset;
  wire  tags_25_clock;
  wire  tags_25_reset;
  wire  tags_26_clock;
  wire  tags_26_reset;
  wire  tags_27_clock;
  wire  tags_27_reset;
  wire  tags_28_clock;
  wire  tags_28_reset;
  wire  tags_29_clock;
  wire  tags_29_reset;
  wire  tags_30_clock;
  wire  tags_30_reset;
  wire  tags_31_clock;
  wire  tags_31_reset;
  wire  tags_32_clock;
  wire  tags_32_reset;
  wire  tags_33_clock;
  wire  tags_33_reset;
  wire  tags_34_clock;
  wire  tags_34_reset;
  wire  tags_35_clock;
  wire  tags_35_reset;
  wire  tags_36_clock;
  wire  tags_36_reset;
  wire  tags_37_clock;
  wire  tags_37_reset;
  wire  tags_38_clock;
  wire  tags_38_reset;
  wire  tags_39_clock;
  wire  tags_39_reset;
  wire  tags_40_clock;
  wire  tags_40_reset;
  wire  tags_41_clock;
  wire  tags_41_reset;
  wire  tags_42_clock;
  wire  tags_42_reset;
  wire  tags_43_clock;
  wire  tags_43_reset;
  wire  tags_44_clock;
  wire  tags_44_reset;
  wire  tags_45_clock;
  wire  tags_45_reset;
  wire  tags_46_clock;
  wire  tags_46_reset;
  wire  tags_47_clock;
  wire  tags_47_reset;
  wire  tags_48_clock;
  wire  tags_48_reset;
  wire  tags_49_clock;
  wire  tags_49_reset;
  wire  tags_50_clock;
  wire  tags_50_reset;
  wire  tags_51_clock;
  wire  tags_51_reset;
  wire  tags_52_clock;
  wire  tags_52_reset;
  wire  tags_53_clock;
  wire  tags_53_reset;
  wire  tags_54_clock;
  wire  tags_54_reset;
  wire  tags_55_clock;
  wire  tags_55_reset;
  wire  tags_56_clock;
  wire  tags_56_reset;
  wire  tags_57_clock;
  wire  tags_57_reset;
  wire  tags_58_clock;
  wire  tags_58_reset;
  wire  tags_59_clock;
  wire  tags_59_reset;
  wire  tags_60_clock;
  wire  tags_60_reset;
  wire  tags_61_clock;
  wire  tags_61_reset;
  wire  tags_62_clock;
  wire  tags_62_reset;
  wire  tags_63_clock;
  wire  tags_63_reset;
  wire  tags_64_clock;
  wire  tags_64_reset;
  wire  tags_65_clock;
  wire  tags_65_reset;
  wire  tags_66_clock;
  wire  tags_66_reset;
  wire  tags_67_clock;
  wire  tags_67_reset;
  wire  tags_68_clock;
  wire  tags_68_reset;
  wire  tags_69_clock;
  wire  tags_69_reset;
  wire  tags_70_clock;
  wire  tags_70_reset;
  wire  tags_71_clock;
  wire  tags_71_reset;
  wire  tags_72_clock;
  wire  tags_72_reset;
  wire  tags_73_clock;
  wire  tags_73_reset;
  wire  tags_74_clock;
  wire  tags_74_reset;
  wire  tags_75_clock;
  wire  tags_75_reset;
  wire  tags_76_clock;
  wire  tags_76_reset;
  wire  tags_77_clock;
  wire  tags_77_reset;
  wire  tags_78_clock;
  wire  tags_78_reset;
  wire  tags_79_clock;
  wire  tags_79_reset;
  wire  tags_80_clock;
  wire  tags_80_reset;
  wire  tags_81_clock;
  wire  tags_81_reset;
  wire  tags_82_clock;
  wire  tags_82_reset;
  wire  tags_83_clock;
  wire  tags_83_reset;
  wire  tags_84_clock;
  wire  tags_84_reset;
  wire  tags_85_clock;
  wire  tags_85_reset;
  wire  tags_86_clock;
  wire  tags_86_reset;
  wire  tags_87_clock;
  wire  tags_87_reset;
  wire  tags_88_clock;
  wire  tags_88_reset;
  wire  tags_89_clock;
  wire  tags_89_reset;
  wire  tags_90_clock;
  wire  tags_90_reset;
  wire  tags_91_clock;
  wire  tags_91_reset;
  wire  tags_92_clock;
  wire  tags_92_reset;
  wire  tags_93_clock;
  wire  tags_93_reset;
  wire  tags_94_clock;
  wire  tags_94_reset;
  wire  tags_95_clock;
  wire  tags_95_reset;
  wire  tags_96_clock;
  wire  tags_96_reset;
  wire  tags_97_clock;
  wire  tags_97_reset;
  wire  tags_98_clock;
  wire  tags_98_reset;
  wire  tags_99_clock;
  wire  tags_99_reset;
  wire  tags_100_clock;
  wire  tags_100_reset;
  wire  tags_101_clock;
  wire  tags_101_reset;
  wire  tags_102_clock;
  wire  tags_102_reset;
  wire  tags_103_clock;
  wire  tags_103_reset;
  wire  tags_104_clock;
  wire  tags_104_reset;
  wire  tags_105_clock;
  wire  tags_105_reset;
  wire  tags_106_clock;
  wire  tags_106_reset;
  wire  tags_107_clock;
  wire  tags_107_reset;
  wire  tags_108_clock;
  wire  tags_108_reset;
  wire  tags_109_clock;
  wire  tags_109_reset;
  wire  tags_110_clock;
  wire  tags_110_reset;
  wire  tags_111_clock;
  wire  tags_111_reset;
  wire  tags_112_clock;
  wire  tags_112_reset;
  wire  tags_113_clock;
  wire  tags_113_reset;
  wire  tags_114_clock;
  wire  tags_114_reset;
  wire  tags_115_clock;
  wire  tags_115_reset;
  wire  tags_116_clock;
  wire  tags_116_reset;
  wire  tags_117_clock;
  wire  tags_117_reset;
  wire  tags_118_clock;
  wire  tags_118_reset;
  wire  tags_119_clock;
  wire  tags_119_reset;
  wire  tags_120_clock;
  wire  tags_120_reset;
  wire  tags_121_clock;
  wire  tags_121_reset;
  wire  tags_122_clock;
  wire  tags_122_reset;
  wire  tags_123_clock;
  wire  tags_123_reset;
  wire  tags_124_clock;
  wire  tags_124_reset;
  wire  tags_125_clock;
  wire  tags_125_reset;
  wire  tags_126_clock;
  wire  tags_126_reset;
  wire  tags_127_clock;
  wire  tags_127_reset;
  wire  tags_128_clock;
  wire  tags_128_reset;
  wire  tags_129_clock;
  wire  tags_129_reset;
  wire  tags_130_clock;
  wire  tags_130_reset;
  wire  tags_131_clock;
  wire  tags_131_reset;
  wire  tags_132_clock;
  wire  tags_132_reset;
  wire  tags_133_clock;
  wire  tags_133_reset;
  wire  tags_134_clock;
  wire  tags_134_reset;
  wire  tags_135_clock;
  wire  tags_135_reset;
  wire  tags_136_clock;
  wire  tags_136_reset;
  wire  tags_137_clock;
  wire  tags_137_reset;
  wire  tags_138_clock;
  wire  tags_138_reset;
  wire  tags_139_clock;
  wire  tags_139_reset;
  wire  tags_140_clock;
  wire  tags_140_reset;
  wire  tags_141_clock;
  wire  tags_141_reset;
  wire  tags_142_clock;
  wire  tags_142_reset;
  wire  tags_143_clock;
  wire  tags_143_reset;
  wire  tags_144_clock;
  wire  tags_144_reset;
  wire  tags_145_clock;
  wire  tags_145_reset;
  wire  tags_146_clock;
  wire  tags_146_reset;
  wire  tags_147_clock;
  wire  tags_147_reset;
  wire  tags_148_clock;
  wire  tags_148_reset;
  wire  tags_149_clock;
  wire  tags_149_reset;
  wire  tags_150_clock;
  wire  tags_150_reset;
  wire  tags_151_clock;
  wire  tags_151_reset;
  wire  tags_152_clock;
  wire  tags_152_reset;
  wire  tags_153_clock;
  wire  tags_153_reset;
  wire  tags_154_clock;
  wire  tags_154_reset;
  wire  tags_155_clock;
  wire  tags_155_reset;
  wire  tags_156_clock;
  wire  tags_156_reset;
  wire  tags_157_clock;
  wire  tags_157_reset;
  wire  tags_158_clock;
  wire  tags_158_reset;
  wire  tags_159_clock;
  wire  tags_159_reset;
  wire  tags_160_clock;
  wire  tags_160_reset;
  wire  tags_161_clock;
  wire  tags_161_reset;
  wire  tags_162_clock;
  wire  tags_162_reset;
  wire  tags_163_clock;
  wire  tags_163_reset;
  wire  tags_164_clock;
  wire  tags_164_reset;
  wire  tags_165_clock;
  wire  tags_165_reset;
  wire  tags_166_clock;
  wire  tags_166_reset;
  wire  tags_167_clock;
  wire  tags_167_reset;
  wire  tags_168_clock;
  wire  tags_168_reset;
  wire  tags_169_clock;
  wire  tags_169_reset;
  wire  tags_170_clock;
  wire  tags_170_reset;
  wire  tags_171_clock;
  wire  tags_171_reset;
  wire  tags_172_clock;
  wire  tags_172_reset;
  wire  tags_173_clock;
  wire  tags_173_reset;
  wire  tags_174_clock;
  wire  tags_174_reset;
  wire  tags_175_clock;
  wire  tags_175_reset;
  wire  tags_176_clock;
  wire  tags_176_reset;
  wire  tags_177_clock;
  wire  tags_177_reset;
  wire  tags_178_clock;
  wire  tags_178_reset;
  wire  tags_179_clock;
  wire  tags_179_reset;
  wire  tags_180_clock;
  wire  tags_180_reset;
  wire  tags_181_clock;
  wire  tags_181_reset;
  wire  tags_182_clock;
  wire  tags_182_reset;
  wire  tags_183_clock;
  wire  tags_183_reset;
  wire  tags_184_clock;
  wire  tags_184_reset;
  wire  tags_185_clock;
  wire  tags_185_reset;
  wire  tags_186_clock;
  wire  tags_186_reset;
  wire  tags_187_clock;
  wire  tags_187_reset;
  wire  tags_188_clock;
  wire  tags_188_reset;
  wire  tags_189_clock;
  wire  tags_189_reset;
  wire  tags_190_clock;
  wire  tags_190_reset;
  wire  tags_191_clock;
  wire  tags_191_reset;
  wire  tags_192_clock;
  wire  tags_192_reset;
  wire  tags_193_clock;
  wire  tags_193_reset;
  wire  tags_194_clock;
  wire  tags_194_reset;
  wire  tags_195_clock;
  wire  tags_195_reset;
  wire  tags_196_clock;
  wire  tags_196_reset;
  wire  tags_197_clock;
  wire  tags_197_reset;
  wire  tags_198_clock;
  wire  tags_198_reset;
  wire  tags_199_clock;
  wire  tags_199_reset;
  wire  tags_200_clock;
  wire  tags_200_reset;
  wire  tags_201_clock;
  wire  tags_201_reset;
  wire  tags_202_clock;
  wire  tags_202_reset;
  wire  tags_203_clock;
  wire  tags_203_reset;
  wire  tags_204_clock;
  wire  tags_204_reset;
  wire  tags_205_clock;
  wire  tags_205_reset;
  wire  tags_206_clock;
  wire  tags_206_reset;
  wire  tags_207_clock;
  wire  tags_207_reset;
  wire  tags_208_clock;
  wire  tags_208_reset;
  wire  tags_209_clock;
  wire  tags_209_reset;
  wire  tags_210_clock;
  wire  tags_210_reset;
  wire  tags_211_clock;
  wire  tags_211_reset;
  wire  tags_212_clock;
  wire  tags_212_reset;
  wire  tags_213_clock;
  wire  tags_213_reset;
  wire  tags_214_clock;
  wire  tags_214_reset;
  wire  tags_215_clock;
  wire  tags_215_reset;
  wire  tags_216_clock;
  wire  tags_216_reset;
  wire  tags_217_clock;
  wire  tags_217_reset;
  wire  tags_218_clock;
  wire  tags_218_reset;
  wire  tags_219_clock;
  wire  tags_219_reset;
  wire  tags_220_clock;
  wire  tags_220_reset;
  wire  tags_221_clock;
  wire  tags_221_reset;
  wire  tags_222_clock;
  wire  tags_222_reset;
  wire  tags_223_clock;
  wire  tags_223_reset;
  wire  tags_224_clock;
  wire  tags_224_reset;
  wire  tags_225_clock;
  wire  tags_225_reset;
  wire  tags_226_clock;
  wire  tags_226_reset;
  wire  tags_227_clock;
  wire  tags_227_reset;
  wire  tags_228_clock;
  wire  tags_228_reset;
  wire  tags_229_clock;
  wire  tags_229_reset;
  wire  tags_230_clock;
  wire  tags_230_reset;
  wire  tags_231_clock;
  wire  tags_231_reset;
  wire  tags_232_clock;
  wire  tags_232_reset;
  wire  tags_233_clock;
  wire  tags_233_reset;
  wire  tags_234_clock;
  wire  tags_234_reset;
  wire  tags_235_clock;
  wire  tags_235_reset;
  wire  tags_236_clock;
  wire  tags_236_reset;
  wire  tags_237_clock;
  wire  tags_237_reset;
  wire  tags_238_clock;
  wire  tags_238_reset;
  wire  tags_239_clock;
  wire  tags_239_reset;
  wire  tags_240_clock;
  wire  tags_240_reset;
  wire  tags_241_clock;
  wire  tags_241_reset;
  wire  tags_242_clock;
  wire  tags_242_reset;
  wire  tags_243_clock;
  wire  tags_243_reset;
  wire  tags_244_clock;
  wire  tags_244_reset;
  wire  tags_245_clock;
  wire  tags_245_reset;
  wire  tags_246_clock;
  wire  tags_246_reset;
  wire  tags_247_clock;
  wire  tags_247_reset;
  wire  tags_248_clock;
  wire  tags_248_reset;
  wire  tags_249_clock;
  wire  tags_249_reset;
  wire  tags_250_clock;
  wire  tags_250_reset;
  wire  tags_251_clock;
  wire  tags_251_reset;
  wire  tags_252_clock;
  wire  tags_252_reset;
  wire  tags_253_clock;
  wire  tags_253_reset;
  wire  tags_254_clock;
  wire  tags_254_reset;
  wire  tags_255_clock;
  wire  tags_255_reset;
  wire  tags_256_clock;
  wire  tags_256_reset;
  wire  tags_257_clock;
  wire  tags_257_reset;
  wire  tags_258_clock;
  wire  tags_258_reset;
  wire  tags_259_clock;
  wire  tags_259_reset;
  wire  tags_260_clock;
  wire  tags_260_reset;
  wire  tags_261_clock;
  wire  tags_261_reset;
  wire  tags_262_clock;
  wire  tags_262_reset;
  wire  tags_263_clock;
  wire  tags_263_reset;
  wire  tags_264_clock;
  wire  tags_264_reset;
  wire  tags_265_clock;
  wire  tags_265_reset;
  wire  tags_266_clock;
  wire  tags_266_reset;
  wire  tags_267_clock;
  wire  tags_267_reset;
  wire  tags_268_clock;
  wire  tags_268_reset;
  wire  tags_269_clock;
  wire  tags_269_reset;
  wire  tags_270_clock;
  wire  tags_270_reset;
  wire  tags_271_clock;
  wire  tags_271_reset;
  wire  tags_272_clock;
  wire  tags_272_reset;
  wire  tags_273_clock;
  wire  tags_273_reset;
  wire  tags_274_clock;
  wire  tags_274_reset;
  wire  tags_275_clock;
  wire  tags_275_reset;
  wire  tags_276_clock;
  wire  tags_276_reset;
  wire  tags_277_clock;
  wire  tags_277_reset;
  wire  tags_278_clock;
  wire  tags_278_reset;
  wire  tags_279_clock;
  wire  tags_279_reset;
  wire  tags_280_clock;
  wire  tags_280_reset;
  wire  tags_281_clock;
  wire  tags_281_reset;
  wire  tags_282_clock;
  wire  tags_282_reset;
  wire  tags_283_clock;
  wire  tags_283_reset;
  wire  tags_284_clock;
  wire  tags_284_reset;
  wire  tags_285_clock;
  wire  tags_285_reset;
  wire  tags_286_clock;
  wire  tags_286_reset;
  wire  tags_287_clock;
  wire  tags_287_reset;
  wire  tags_288_clock;
  wire  tags_288_reset;
  wire  tags_289_clock;
  wire  tags_289_reset;
  wire  tags_290_clock;
  wire  tags_290_reset;
  wire  tags_291_clock;
  wire  tags_291_reset;
  wire  tags_292_clock;
  wire  tags_292_reset;
  wire  tags_293_clock;
  wire  tags_293_reset;
  wire  tags_294_clock;
  wire  tags_294_reset;
  wire  tags_295_clock;
  wire  tags_295_reset;
  wire  tags_296_clock;
  wire  tags_296_reset;
  wire  tags_297_clock;
  wire  tags_297_reset;
  wire  tags_298_clock;
  wire  tags_298_reset;
  wire  tags_299_clock;
  wire  tags_299_reset;
  wire  tags_300_clock;
  wire  tags_300_reset;
  wire  tags_301_clock;
  wire  tags_301_reset;
  wire  tags_302_clock;
  wire  tags_302_reset;
  wire  tags_303_clock;
  wire  tags_303_reset;
  wire  tags_304_clock;
  wire  tags_304_reset;
  wire  tags_305_clock;
  wire  tags_305_reset;
  wire  tags_306_clock;
  wire  tags_306_reset;
  wire  tags_307_clock;
  wire  tags_307_reset;
  wire  tags_308_clock;
  wire  tags_308_reset;
  wire  tags_309_clock;
  wire  tags_309_reset;
  wire  tags_310_clock;
  wire  tags_310_reset;
  wire  tags_311_clock;
  wire  tags_311_reset;
  wire  tags_312_clock;
  wire  tags_312_reset;
  wire  tags_313_clock;
  wire  tags_313_reset;
  wire  tags_314_clock;
  wire  tags_314_reset;
  wire  tags_315_clock;
  wire  tags_315_reset;
  wire  tags_316_clock;
  wire  tags_316_reset;
  wire  tags_317_clock;
  wire  tags_317_reset;
  wire  tags_318_clock;
  wire  tags_318_reset;
  wire  tags_319_clock;
  wire  tags_319_reset;
  wire  tags_320_clock;
  wire  tags_320_reset;
  wire  tags_321_clock;
  wire  tags_321_reset;
  wire  tags_322_clock;
  wire  tags_322_reset;
  wire  tags_323_clock;
  wire  tags_323_reset;
  wire  tags_324_clock;
  wire  tags_324_reset;
  wire  tags_325_clock;
  wire  tags_325_reset;
  wire  tags_326_clock;
  wire  tags_326_reset;
  wire  tags_327_clock;
  wire  tags_327_reset;
  wire  tags_328_clock;
  wire  tags_328_reset;
  wire  tags_329_clock;
  wire  tags_329_reset;
  wire  tags_330_clock;
  wire  tags_330_reset;
  wire  tags_331_clock;
  wire  tags_331_reset;
  wire  tags_332_clock;
  wire  tags_332_reset;
  wire  tags_333_clock;
  wire  tags_333_reset;
  wire  tags_334_clock;
  wire  tags_334_reset;
  wire  tags_335_clock;
  wire  tags_335_reset;
  wire  tags_336_clock;
  wire  tags_336_reset;
  wire  tags_337_clock;
  wire  tags_337_reset;
  wire  tags_338_clock;
  wire  tags_338_reset;
  wire  tags_339_clock;
  wire  tags_339_reset;
  wire  tags_340_clock;
  wire  tags_340_reset;
  wire  tags_341_clock;
  wire  tags_341_reset;
  wire  tags_342_clock;
  wire  tags_342_reset;
  wire  tags_343_clock;
  wire  tags_343_reset;
  wire  tags_344_clock;
  wire  tags_344_reset;
  wire  tags_345_clock;
  wire  tags_345_reset;
  wire  tags_346_clock;
  wire  tags_346_reset;
  wire  tags_347_clock;
  wire  tags_347_reset;
  wire  tags_348_clock;
  wire  tags_348_reset;
  wire  tags_349_clock;
  wire  tags_349_reset;
  wire  tags_350_clock;
  wire  tags_350_reset;
  wire  tags_351_clock;
  wire  tags_351_reset;
  wire  tags_352_clock;
  wire  tags_352_reset;
  wire  tags_353_clock;
  wire  tags_353_reset;
  wire  tags_354_clock;
  wire  tags_354_reset;
  wire  tags_355_clock;
  wire  tags_355_reset;
  wire  tags_356_clock;
  wire  tags_356_reset;
  wire  tags_357_clock;
  wire  tags_357_reset;
  wire  tags_358_clock;
  wire  tags_358_reset;
  wire  tags_359_clock;
  wire  tags_359_reset;
  wire  tags_360_clock;
  wire  tags_360_reset;
  wire  tags_361_clock;
  wire  tags_361_reset;
  wire  tags_362_clock;
  wire  tags_362_reset;
  wire  tags_363_clock;
  wire  tags_363_reset;
  wire  tags_364_clock;
  wire  tags_364_reset;
  wire  tags_365_clock;
  wire  tags_365_reset;
  wire  tags_366_clock;
  wire  tags_366_reset;
  wire  tags_367_clock;
  wire  tags_367_reset;
  wire  tags_368_clock;
  wire  tags_368_reset;
  wire  tags_369_clock;
  wire  tags_369_reset;
  wire  tags_370_clock;
  wire  tags_370_reset;
  wire  tags_371_clock;
  wire  tags_371_reset;
  wire  tags_372_clock;
  wire  tags_372_reset;
  wire  tags_373_clock;
  wire  tags_373_reset;
  wire  tags_374_clock;
  wire  tags_374_reset;
  wire  tags_375_clock;
  wire  tags_375_reset;
  wire  tags_376_clock;
  wire  tags_376_reset;
  wire  tags_377_clock;
  wire  tags_377_reset;
  wire  tags_378_clock;
  wire  tags_378_reset;
  wire  tags_379_clock;
  wire  tags_379_reset;
  wire  tags_380_clock;
  wire  tags_380_reset;
  wire  tags_381_clock;
  wire  tags_381_reset;
  wire  tags_382_clock;
  wire  tags_382_reset;
  wire  tags_383_clock;
  wire  tags_383_reset;
  wire  tags_384_clock;
  wire  tags_384_reset;
  wire  tags_385_clock;
  wire  tags_385_reset;
  wire  tags_386_clock;
  wire  tags_386_reset;
  wire  tags_387_clock;
  wire  tags_387_reset;
  wire  tags_388_clock;
  wire  tags_388_reset;
  wire  tags_389_clock;
  wire  tags_389_reset;
  wire  tags_390_clock;
  wire  tags_390_reset;
  wire  tags_391_clock;
  wire  tags_391_reset;
  wire  tags_392_clock;
  wire  tags_392_reset;
  wire  tags_393_clock;
  wire  tags_393_reset;
  wire  tags_394_clock;
  wire  tags_394_reset;
  wire  tags_395_clock;
  wire  tags_395_reset;
  wire  tags_396_clock;
  wire  tags_396_reset;
  wire  tags_397_clock;
  wire  tags_397_reset;
  wire  tags_398_clock;
  wire  tags_398_reset;
  wire  tags_399_clock;
  wire  tags_399_reset;
  wire  tags_400_clock;
  wire  tags_400_reset;
  wire  tags_401_clock;
  wire  tags_401_reset;
  wire  tags_402_clock;
  wire  tags_402_reset;
  wire  tags_403_clock;
  wire  tags_403_reset;
  wire  tags_404_clock;
  wire  tags_404_reset;
  wire  tags_405_clock;
  wire  tags_405_reset;
  wire  tags_406_clock;
  wire  tags_406_reset;
  wire  tags_407_clock;
  wire  tags_407_reset;
  wire  tags_408_clock;
  wire  tags_408_reset;
  wire  tags_409_clock;
  wire  tags_409_reset;
  wire  tags_410_clock;
  wire  tags_410_reset;
  wire  tags_411_clock;
  wire  tags_411_reset;
  wire  tags_412_clock;
  wire  tags_412_reset;
  wire  tags_413_clock;
  wire  tags_413_reset;
  wire  tags_414_clock;
  wire  tags_414_reset;
  wire  tags_415_clock;
  wire  tags_415_reset;
  wire  tags_416_clock;
  wire  tags_416_reset;
  wire  tags_417_clock;
  wire  tags_417_reset;
  wire  tags_418_clock;
  wire  tags_418_reset;
  wire  tags_419_clock;
  wire  tags_419_reset;
  wire  tags_420_clock;
  wire  tags_420_reset;
  wire  tags_421_clock;
  wire  tags_421_reset;
  wire  tags_422_clock;
  wire  tags_422_reset;
  wire  tags_423_clock;
  wire  tags_423_reset;
  wire  tags_424_clock;
  wire  tags_424_reset;
  wire  tags_425_clock;
  wire  tags_425_reset;
  wire  tags_426_clock;
  wire  tags_426_reset;
  wire  tags_427_clock;
  wire  tags_427_reset;
  wire  tags_428_clock;
  wire  tags_428_reset;
  wire  tags_429_clock;
  wire  tags_429_reset;
  wire  tags_430_clock;
  wire  tags_430_reset;
  wire  tags_431_clock;
  wire  tags_431_reset;
  wire  tags_432_clock;
  wire  tags_432_reset;
  wire  tags_433_clock;
  wire  tags_433_reset;
  wire  tags_434_clock;
  wire  tags_434_reset;
  wire  tags_435_clock;
  wire  tags_435_reset;
  wire  tags_436_clock;
  wire  tags_436_reset;
  wire  tags_437_clock;
  wire  tags_437_reset;
  wire  tags_438_clock;
  wire  tags_438_reset;
  wire  tags_439_clock;
  wire  tags_439_reset;
  wire  tags_440_clock;
  wire  tags_440_reset;
  wire  tags_441_clock;
  wire  tags_441_reset;
  wire  tags_442_clock;
  wire  tags_442_reset;
  wire  tags_443_clock;
  wire  tags_443_reset;
  wire  tags_444_clock;
  wire  tags_444_reset;
  wire  tags_445_clock;
  wire  tags_445_reset;
  wire  tags_446_clock;
  wire  tags_446_reset;
  wire  tags_447_clock;
  wire  tags_447_reset;
  wire  tags_448_clock;
  wire  tags_448_reset;
  wire  tags_449_clock;
  wire  tags_449_reset;
  wire  tags_450_clock;
  wire  tags_450_reset;
  wire  tags_451_clock;
  wire  tags_451_reset;
  wire  tags_452_clock;
  wire  tags_452_reset;
  wire  tags_453_clock;
  wire  tags_453_reset;
  wire  tags_454_clock;
  wire  tags_454_reset;
  wire  tags_455_clock;
  wire  tags_455_reset;
  wire  tags_456_clock;
  wire  tags_456_reset;
  wire  tags_457_clock;
  wire  tags_457_reset;
  wire  tags_458_clock;
  wire  tags_458_reset;
  wire  tags_459_clock;
  wire  tags_459_reset;
  wire  tags_460_clock;
  wire  tags_460_reset;
  wire  tags_461_clock;
  wire  tags_461_reset;
  wire  tags_462_clock;
  wire  tags_462_reset;
  wire  tags_463_clock;
  wire  tags_463_reset;
  wire  tags_464_clock;
  wire  tags_464_reset;
  wire  tags_465_clock;
  wire  tags_465_reset;
  wire  tags_466_clock;
  wire  tags_466_reset;
  wire  tags_467_clock;
  wire  tags_467_reset;
  wire  tags_468_clock;
  wire  tags_468_reset;
  wire  tags_469_clock;
  wire  tags_469_reset;
  wire  tags_470_clock;
  wire  tags_470_reset;
  wire  tags_471_clock;
  wire  tags_471_reset;
  wire  tags_472_clock;
  wire  tags_472_reset;
  wire  tags_473_clock;
  wire  tags_473_reset;
  wire  tags_474_clock;
  wire  tags_474_reset;
  wire  tags_475_clock;
  wire  tags_475_reset;
  wire  tags_476_clock;
  wire  tags_476_reset;
  wire  tags_477_clock;
  wire  tags_477_reset;
  wire  tags_478_clock;
  wire  tags_478_reset;
  wire  tags_479_clock;
  wire  tags_479_reset;
  wire  tags_480_clock;
  wire  tags_480_reset;
  wire  tags_481_clock;
  wire  tags_481_reset;
  wire  tags_482_clock;
  wire  tags_482_reset;
  wire  tags_483_clock;
  wire  tags_483_reset;
  wire  tags_484_clock;
  wire  tags_484_reset;
  wire  tags_485_clock;
  wire  tags_485_reset;
  wire  tags_486_clock;
  wire  tags_486_reset;
  wire  tags_487_clock;
  wire  tags_487_reset;
  wire  tags_488_clock;
  wire  tags_488_reset;
  wire  tags_489_clock;
  wire  tags_489_reset;
  wire  tags_490_clock;
  wire  tags_490_reset;
  wire  tags_491_clock;
  wire  tags_491_reset;
  wire  tags_492_clock;
  wire  tags_492_reset;
  wire  tags_493_clock;
  wire  tags_493_reset;
  wire  tags_494_clock;
  wire  tags_494_reset;
  wire  tags_495_clock;
  wire  tags_495_reset;
  wire  tags_496_clock;
  wire  tags_496_reset;
  wire  tags_497_clock;
  wire  tags_497_reset;
  wire  tags_498_clock;
  wire  tags_498_reset;
  wire  tags_499_clock;
  wire  tags_499_reset;
  wire  tags_500_clock;
  wire  tags_500_reset;
  wire  tags_501_clock;
  wire  tags_501_reset;
  wire  tags_502_clock;
  wire  tags_502_reset;
  wire  tags_503_clock;
  wire  tags_503_reset;
  wire  tags_504_clock;
  wire  tags_504_reset;
  wire  tags_505_clock;
  wire  tags_505_reset;
  wire  tags_506_clock;
  wire  tags_506_reset;
  wire  tags_507_clock;
  wire  tags_507_reset;
  wire  tags_508_clock;
  wire  tags_508_reset;
  wire  tags_509_clock;
  wire  tags_509_reset;
  wire  tags_510_clock;
  wire  tags_510_reset;
  wire  tags_511_clock;
  wire  tags_511_reset;
  wire  metadata_clock;
  wire [7:0] metadata_io_wdata_0;
  wire [7:0] metadata_io_wdata_1;
  wire [7:0] metadata_io_wdata_2;
  wire [7:0] metadata_io_wdata_3;
  wire [7:0] metadata_io_wdata_4;
  wire [7:0] metadata_io_wdata_5;
  wire [7:0] metadata_io_wdata_6;
  wire [7:0] metadata_io_wdata_7;
  wire [7:0] metadata_io_wdata_8;
  wire [7:0] metadata_io_wdata_9;
  wire [7:0] metadata_io_wdata_10;
  wire [7:0] metadata_io_wdata_11;
  wire [7:0] metadata_io_wdata_12;
  wire [7:0] metadata_io_wdata_13;
  wire [7:0] metadata_io_wdata_14;
  wire [7:0] metadata_io_wdata_15;
  wire [7:0] metadata_io_rdata_0;
  wire [7:0] metadata_io_rdata_1;
  wire [7:0] metadata_io_rdata_2;
  wire [7:0] metadata_io_rdata_3;
  wire [7:0] metadata_io_rdata_4;
  wire [7:0] metadata_io_rdata_5;
  wire [7:0] metadata_io_rdata_6;
  wire [7:0] metadata_io_rdata_7;
  wire [7:0] metadata_io_rdata_8;
  wire [7:0] metadata_io_rdata_9;
  wire [7:0] metadata_io_rdata_10;
  wire [7:0] metadata_io_rdata_11;
  wire [7:0] metadata_io_rdata_12;
  wire [7:0] metadata_io_rdata_13;
  wire [7:0] metadata_io_rdata_14;
  wire [7:0] metadata_io_rdata_15;
  wire [3:0] woffset;
  wire [3:0] _T_19089;
  wire [7:0] md_0;
  wire [7:0] md_1;
  wire [7:0] md_2;
  wire [7:0] md_3;
  wire [7:0] md_4;
  wire [7:0] md_5;
  wire [7:0] md_6;
  wire [7:0] md_7;
  wire [7:0] md_8;
  wire [7:0] md_9;
  wire [7:0] md_10;
  wire [7:0] md_11;
  wire [7:0] md_12;
  wire [7:0] md_13;
  wire [7:0] md_14;
  wire [7:0] md_15;
  wire [4:0] _T_19127;
  wire [7:0] _GEN_0;
  wire [7:0] _GEN_2;
  wire [7:0] _GEN_3;
  wire [7:0] _GEN_4;
  wire [7:0] _GEN_5;
  wire [7:0] _GEN_6;
  wire [7:0] _GEN_7;
  wire [7:0] _GEN_8;
  wire [7:0] _GEN_9;
  wire [7:0] _GEN_10;
  wire [7:0] _GEN_11;
  wire [7:0] _GEN_12;
  wire [7:0] _GEN_13;
  wire [7:0] _GEN_14;
  wire [7:0] _GEN_15;
  wire [7:0] _GEN_16;
  wire [7:0] _GEN_17;
  FF_9 valid_0 (
    .clock(valid_0_clock),
    .reset(valid_0_reset),
    .io_in(valid_0_io_in),
    .io_out(valid_0_io_out),
    .io_enable(valid_0_io_enable)
  );
  FF_9 valid_1 (
    .clock(valid_1_clock),
    .reset(valid_1_reset),
    .io_in(valid_1_io_in),
    .io_out(valid_1_io_out),
    .io_enable(valid_1_io_enable)
  );
  FF_9 valid_2 (
    .clock(valid_2_clock),
    .reset(valid_2_reset),
    .io_in(valid_2_io_in),
    .io_out(valid_2_io_out),
    .io_enable(valid_2_io_enable)
  );
  FF_9 valid_3 (
    .clock(valid_3_clock),
    .reset(valid_3_reset),
    .io_in(valid_3_io_in),
    .io_out(valid_3_io_out),
    .io_enable(valid_3_io_enable)
  );
  FF_9 valid_4 (
    .clock(valid_4_clock),
    .reset(valid_4_reset),
    .io_in(valid_4_io_in),
    .io_out(valid_4_io_out),
    .io_enable(valid_4_io_enable)
  );
  FF_9 valid_5 (
    .clock(valid_5_clock),
    .reset(valid_5_reset),
    .io_in(valid_5_io_in),
    .io_out(valid_5_io_out),
    .io_enable(valid_5_io_enable)
  );
  FF_9 valid_6 (
    .clock(valid_6_clock),
    .reset(valid_6_reset),
    .io_in(valid_6_io_in),
    .io_out(valid_6_io_out),
    .io_enable(valid_6_io_enable)
  );
  FF_9 valid_7 (
    .clock(valid_7_clock),
    .reset(valid_7_reset),
    .io_in(valid_7_io_in),
    .io_out(valid_7_io_out),
    .io_enable(valid_7_io_enable)
  );
  FF_9 valid_8 (
    .clock(valid_8_clock),
    .reset(valid_8_reset),
    .io_in(valid_8_io_in),
    .io_out(valid_8_io_out),
    .io_enable(valid_8_io_enable)
  );
  FF_9 valid_9 (
    .clock(valid_9_clock),
    .reset(valid_9_reset),
    .io_in(valid_9_io_in),
    .io_out(valid_9_io_out),
    .io_enable(valid_9_io_enable)
  );
  FF_9 valid_10 (
    .clock(valid_10_clock),
    .reset(valid_10_reset),
    .io_in(valid_10_io_in),
    .io_out(valid_10_io_out),
    .io_enable(valid_10_io_enable)
  );
  FF_9 valid_11 (
    .clock(valid_11_clock),
    .reset(valid_11_reset),
    .io_in(valid_11_io_in),
    .io_out(valid_11_io_out),
    .io_enable(valid_11_io_enable)
  );
  FF_9 valid_12 (
    .clock(valid_12_clock),
    .reset(valid_12_reset),
    .io_in(valid_12_io_in),
    .io_out(valid_12_io_out),
    .io_enable(valid_12_io_enable)
  );
  FF_9 valid_13 (
    .clock(valid_13_clock),
    .reset(valid_13_reset),
    .io_in(valid_13_io_in),
    .io_out(valid_13_io_out),
    .io_enable(valid_13_io_enable)
  );
  FF_9 valid_14 (
    .clock(valid_14_clock),
    .reset(valid_14_reset),
    .io_in(valid_14_io_in),
    .io_out(valid_14_io_out),
    .io_enable(valid_14_io_enable)
  );
  FF_9 valid_15 (
    .clock(valid_15_clock),
    .reset(valid_15_reset),
    .io_in(valid_15_io_in),
    .io_out(valid_15_io_out),
    .io_enable(valid_15_io_enable)
  );
  FF_9 valid_16 (
    .clock(valid_16_clock),
    .reset(valid_16_reset),
    .io_in(valid_16_io_in),
    .io_out(valid_16_io_out),
    .io_enable(valid_16_io_enable)
  );
  FF_9 valid_17 (
    .clock(valid_17_clock),
    .reset(valid_17_reset),
    .io_in(valid_17_io_in),
    .io_out(valid_17_io_out),
    .io_enable(valid_17_io_enable)
  );
  FF_9 valid_18 (
    .clock(valid_18_clock),
    .reset(valid_18_reset),
    .io_in(valid_18_io_in),
    .io_out(valid_18_io_out),
    .io_enable(valid_18_io_enable)
  );
  FF_9 valid_19 (
    .clock(valid_19_clock),
    .reset(valid_19_reset),
    .io_in(valid_19_io_in),
    .io_out(valid_19_io_out),
    .io_enable(valid_19_io_enable)
  );
  FF_9 valid_20 (
    .clock(valid_20_clock),
    .reset(valid_20_reset),
    .io_in(valid_20_io_in),
    .io_out(valid_20_io_out),
    .io_enable(valid_20_io_enable)
  );
  FF_9 valid_21 (
    .clock(valid_21_clock),
    .reset(valid_21_reset),
    .io_in(valid_21_io_in),
    .io_out(valid_21_io_out),
    .io_enable(valid_21_io_enable)
  );
  FF_9 valid_22 (
    .clock(valid_22_clock),
    .reset(valid_22_reset),
    .io_in(valid_22_io_in),
    .io_out(valid_22_io_out),
    .io_enable(valid_22_io_enable)
  );
  FF_9 valid_23 (
    .clock(valid_23_clock),
    .reset(valid_23_reset),
    .io_in(valid_23_io_in),
    .io_out(valid_23_io_out),
    .io_enable(valid_23_io_enable)
  );
  FF_9 valid_24 (
    .clock(valid_24_clock),
    .reset(valid_24_reset),
    .io_in(valid_24_io_in),
    .io_out(valid_24_io_out),
    .io_enable(valid_24_io_enable)
  );
  FF_9 valid_25 (
    .clock(valid_25_clock),
    .reset(valid_25_reset),
    .io_in(valid_25_io_in),
    .io_out(valid_25_io_out),
    .io_enable(valid_25_io_enable)
  );
  FF_9 valid_26 (
    .clock(valid_26_clock),
    .reset(valid_26_reset),
    .io_in(valid_26_io_in),
    .io_out(valid_26_io_out),
    .io_enable(valid_26_io_enable)
  );
  FF_9 valid_27 (
    .clock(valid_27_clock),
    .reset(valid_27_reset),
    .io_in(valid_27_io_in),
    .io_out(valid_27_io_out),
    .io_enable(valid_27_io_enable)
  );
  FF_9 valid_28 (
    .clock(valid_28_clock),
    .reset(valid_28_reset),
    .io_in(valid_28_io_in),
    .io_out(valid_28_io_out),
    .io_enable(valid_28_io_enable)
  );
  FF_9 valid_29 (
    .clock(valid_29_clock),
    .reset(valid_29_reset),
    .io_in(valid_29_io_in),
    .io_out(valid_29_io_out),
    .io_enable(valid_29_io_enable)
  );
  FF_9 valid_30 (
    .clock(valid_30_clock),
    .reset(valid_30_reset),
    .io_in(valid_30_io_in),
    .io_out(valid_30_io_out),
    .io_enable(valid_30_io_enable)
  );
  FF_9 valid_31 (
    .clock(valid_31_clock),
    .reset(valid_31_reset),
    .io_in(valid_31_io_in),
    .io_out(valid_31_io_out),
    .io_enable(valid_31_io_enable)
  );
  FF_9 valid_32 (
    .clock(valid_32_clock),
    .reset(valid_32_reset),
    .io_in(valid_32_io_in),
    .io_out(valid_32_io_out),
    .io_enable(valid_32_io_enable)
  );
  FF_9 valid_33 (
    .clock(valid_33_clock),
    .reset(valid_33_reset),
    .io_in(valid_33_io_in),
    .io_out(valid_33_io_out),
    .io_enable(valid_33_io_enable)
  );
  FF_9 valid_34 (
    .clock(valid_34_clock),
    .reset(valid_34_reset),
    .io_in(valid_34_io_in),
    .io_out(valid_34_io_out),
    .io_enable(valid_34_io_enable)
  );
  FF_9 valid_35 (
    .clock(valid_35_clock),
    .reset(valid_35_reset),
    .io_in(valid_35_io_in),
    .io_out(valid_35_io_out),
    .io_enable(valid_35_io_enable)
  );
  FF_9 valid_36 (
    .clock(valid_36_clock),
    .reset(valid_36_reset),
    .io_in(valid_36_io_in),
    .io_out(valid_36_io_out),
    .io_enable(valid_36_io_enable)
  );
  FF_9 valid_37 (
    .clock(valid_37_clock),
    .reset(valid_37_reset),
    .io_in(valid_37_io_in),
    .io_out(valid_37_io_out),
    .io_enable(valid_37_io_enable)
  );
  FF_9 valid_38 (
    .clock(valid_38_clock),
    .reset(valid_38_reset),
    .io_in(valid_38_io_in),
    .io_out(valid_38_io_out),
    .io_enable(valid_38_io_enable)
  );
  FF_9 valid_39 (
    .clock(valid_39_clock),
    .reset(valid_39_reset),
    .io_in(valid_39_io_in),
    .io_out(valid_39_io_out),
    .io_enable(valid_39_io_enable)
  );
  FF_9 valid_40 (
    .clock(valid_40_clock),
    .reset(valid_40_reset),
    .io_in(valid_40_io_in),
    .io_out(valid_40_io_out),
    .io_enable(valid_40_io_enable)
  );
  FF_9 valid_41 (
    .clock(valid_41_clock),
    .reset(valid_41_reset),
    .io_in(valid_41_io_in),
    .io_out(valid_41_io_out),
    .io_enable(valid_41_io_enable)
  );
  FF_9 valid_42 (
    .clock(valid_42_clock),
    .reset(valid_42_reset),
    .io_in(valid_42_io_in),
    .io_out(valid_42_io_out),
    .io_enable(valid_42_io_enable)
  );
  FF_9 valid_43 (
    .clock(valid_43_clock),
    .reset(valid_43_reset),
    .io_in(valid_43_io_in),
    .io_out(valid_43_io_out),
    .io_enable(valid_43_io_enable)
  );
  FF_9 valid_44 (
    .clock(valid_44_clock),
    .reset(valid_44_reset),
    .io_in(valid_44_io_in),
    .io_out(valid_44_io_out),
    .io_enable(valid_44_io_enable)
  );
  FF_9 valid_45 (
    .clock(valid_45_clock),
    .reset(valid_45_reset),
    .io_in(valid_45_io_in),
    .io_out(valid_45_io_out),
    .io_enable(valid_45_io_enable)
  );
  FF_9 valid_46 (
    .clock(valid_46_clock),
    .reset(valid_46_reset),
    .io_in(valid_46_io_in),
    .io_out(valid_46_io_out),
    .io_enable(valid_46_io_enable)
  );
  FF_9 valid_47 (
    .clock(valid_47_clock),
    .reset(valid_47_reset),
    .io_in(valid_47_io_in),
    .io_out(valid_47_io_out),
    .io_enable(valid_47_io_enable)
  );
  FF_9 valid_48 (
    .clock(valid_48_clock),
    .reset(valid_48_reset),
    .io_in(valid_48_io_in),
    .io_out(valid_48_io_out),
    .io_enable(valid_48_io_enable)
  );
  FF_9 valid_49 (
    .clock(valid_49_clock),
    .reset(valid_49_reset),
    .io_in(valid_49_io_in),
    .io_out(valid_49_io_out),
    .io_enable(valid_49_io_enable)
  );
  FF_9 valid_50 (
    .clock(valid_50_clock),
    .reset(valid_50_reset),
    .io_in(valid_50_io_in),
    .io_out(valid_50_io_out),
    .io_enable(valid_50_io_enable)
  );
  FF_9 valid_51 (
    .clock(valid_51_clock),
    .reset(valid_51_reset),
    .io_in(valid_51_io_in),
    .io_out(valid_51_io_out),
    .io_enable(valid_51_io_enable)
  );
  FF_9 valid_52 (
    .clock(valid_52_clock),
    .reset(valid_52_reset),
    .io_in(valid_52_io_in),
    .io_out(valid_52_io_out),
    .io_enable(valid_52_io_enable)
  );
  FF_9 valid_53 (
    .clock(valid_53_clock),
    .reset(valid_53_reset),
    .io_in(valid_53_io_in),
    .io_out(valid_53_io_out),
    .io_enable(valid_53_io_enable)
  );
  FF_9 valid_54 (
    .clock(valid_54_clock),
    .reset(valid_54_reset),
    .io_in(valid_54_io_in),
    .io_out(valid_54_io_out),
    .io_enable(valid_54_io_enable)
  );
  FF_9 valid_55 (
    .clock(valid_55_clock),
    .reset(valid_55_reset),
    .io_in(valid_55_io_in),
    .io_out(valid_55_io_out),
    .io_enable(valid_55_io_enable)
  );
  FF_9 valid_56 (
    .clock(valid_56_clock),
    .reset(valid_56_reset),
    .io_in(valid_56_io_in),
    .io_out(valid_56_io_out),
    .io_enable(valid_56_io_enable)
  );
  FF_9 valid_57 (
    .clock(valid_57_clock),
    .reset(valid_57_reset),
    .io_in(valid_57_io_in),
    .io_out(valid_57_io_out),
    .io_enable(valid_57_io_enable)
  );
  FF_9 valid_58 (
    .clock(valid_58_clock),
    .reset(valid_58_reset),
    .io_in(valid_58_io_in),
    .io_out(valid_58_io_out),
    .io_enable(valid_58_io_enable)
  );
  FF_9 valid_59 (
    .clock(valid_59_clock),
    .reset(valid_59_reset),
    .io_in(valid_59_io_in),
    .io_out(valid_59_io_out),
    .io_enable(valid_59_io_enable)
  );
  FF_9 valid_60 (
    .clock(valid_60_clock),
    .reset(valid_60_reset),
    .io_in(valid_60_io_in),
    .io_out(valid_60_io_out),
    .io_enable(valid_60_io_enable)
  );
  FF_9 valid_61 (
    .clock(valid_61_clock),
    .reset(valid_61_reset),
    .io_in(valid_61_io_in),
    .io_out(valid_61_io_out),
    .io_enable(valid_61_io_enable)
  );
  FF_9 valid_62 (
    .clock(valid_62_clock),
    .reset(valid_62_reset),
    .io_in(valid_62_io_in),
    .io_out(valid_62_io_out),
    .io_enable(valid_62_io_enable)
  );
  FF_9 valid_63 (
    .clock(valid_63_clock),
    .reset(valid_63_reset),
    .io_in(valid_63_io_in),
    .io_out(valid_63_io_out),
    .io_enable(valid_63_io_enable)
  );
  FF_9 valid_64 (
    .clock(valid_64_clock),
    .reset(valid_64_reset),
    .io_in(valid_64_io_in),
    .io_out(valid_64_io_out),
    .io_enable(valid_64_io_enable)
  );
  FF_9 valid_65 (
    .clock(valid_65_clock),
    .reset(valid_65_reset),
    .io_in(valid_65_io_in),
    .io_out(valid_65_io_out),
    .io_enable(valid_65_io_enable)
  );
  FF_9 valid_66 (
    .clock(valid_66_clock),
    .reset(valid_66_reset),
    .io_in(valid_66_io_in),
    .io_out(valid_66_io_out),
    .io_enable(valid_66_io_enable)
  );
  FF_9 valid_67 (
    .clock(valid_67_clock),
    .reset(valid_67_reset),
    .io_in(valid_67_io_in),
    .io_out(valid_67_io_out),
    .io_enable(valid_67_io_enable)
  );
  FF_9 valid_68 (
    .clock(valid_68_clock),
    .reset(valid_68_reset),
    .io_in(valid_68_io_in),
    .io_out(valid_68_io_out),
    .io_enable(valid_68_io_enable)
  );
  FF_9 valid_69 (
    .clock(valid_69_clock),
    .reset(valid_69_reset),
    .io_in(valid_69_io_in),
    .io_out(valid_69_io_out),
    .io_enable(valid_69_io_enable)
  );
  FF_9 valid_70 (
    .clock(valid_70_clock),
    .reset(valid_70_reset),
    .io_in(valid_70_io_in),
    .io_out(valid_70_io_out),
    .io_enable(valid_70_io_enable)
  );
  FF_9 valid_71 (
    .clock(valid_71_clock),
    .reset(valid_71_reset),
    .io_in(valid_71_io_in),
    .io_out(valid_71_io_out),
    .io_enable(valid_71_io_enable)
  );
  FF_9 valid_72 (
    .clock(valid_72_clock),
    .reset(valid_72_reset),
    .io_in(valid_72_io_in),
    .io_out(valid_72_io_out),
    .io_enable(valid_72_io_enable)
  );
  FF_9 valid_73 (
    .clock(valid_73_clock),
    .reset(valid_73_reset),
    .io_in(valid_73_io_in),
    .io_out(valid_73_io_out),
    .io_enable(valid_73_io_enable)
  );
  FF_9 valid_74 (
    .clock(valid_74_clock),
    .reset(valid_74_reset),
    .io_in(valid_74_io_in),
    .io_out(valid_74_io_out),
    .io_enable(valid_74_io_enable)
  );
  FF_9 valid_75 (
    .clock(valid_75_clock),
    .reset(valid_75_reset),
    .io_in(valid_75_io_in),
    .io_out(valid_75_io_out),
    .io_enable(valid_75_io_enable)
  );
  FF_9 valid_76 (
    .clock(valid_76_clock),
    .reset(valid_76_reset),
    .io_in(valid_76_io_in),
    .io_out(valid_76_io_out),
    .io_enable(valid_76_io_enable)
  );
  FF_9 valid_77 (
    .clock(valid_77_clock),
    .reset(valid_77_reset),
    .io_in(valid_77_io_in),
    .io_out(valid_77_io_out),
    .io_enable(valid_77_io_enable)
  );
  FF_9 valid_78 (
    .clock(valid_78_clock),
    .reset(valid_78_reset),
    .io_in(valid_78_io_in),
    .io_out(valid_78_io_out),
    .io_enable(valid_78_io_enable)
  );
  FF_9 valid_79 (
    .clock(valid_79_clock),
    .reset(valid_79_reset),
    .io_in(valid_79_io_in),
    .io_out(valid_79_io_out),
    .io_enable(valid_79_io_enable)
  );
  FF_9 valid_80 (
    .clock(valid_80_clock),
    .reset(valid_80_reset),
    .io_in(valid_80_io_in),
    .io_out(valid_80_io_out),
    .io_enable(valid_80_io_enable)
  );
  FF_9 valid_81 (
    .clock(valid_81_clock),
    .reset(valid_81_reset),
    .io_in(valid_81_io_in),
    .io_out(valid_81_io_out),
    .io_enable(valid_81_io_enable)
  );
  FF_9 valid_82 (
    .clock(valid_82_clock),
    .reset(valid_82_reset),
    .io_in(valid_82_io_in),
    .io_out(valid_82_io_out),
    .io_enable(valid_82_io_enable)
  );
  FF_9 valid_83 (
    .clock(valid_83_clock),
    .reset(valid_83_reset),
    .io_in(valid_83_io_in),
    .io_out(valid_83_io_out),
    .io_enable(valid_83_io_enable)
  );
  FF_9 valid_84 (
    .clock(valid_84_clock),
    .reset(valid_84_reset),
    .io_in(valid_84_io_in),
    .io_out(valid_84_io_out),
    .io_enable(valid_84_io_enable)
  );
  FF_9 valid_85 (
    .clock(valid_85_clock),
    .reset(valid_85_reset),
    .io_in(valid_85_io_in),
    .io_out(valid_85_io_out),
    .io_enable(valid_85_io_enable)
  );
  FF_9 valid_86 (
    .clock(valid_86_clock),
    .reset(valid_86_reset),
    .io_in(valid_86_io_in),
    .io_out(valid_86_io_out),
    .io_enable(valid_86_io_enable)
  );
  FF_9 valid_87 (
    .clock(valid_87_clock),
    .reset(valid_87_reset),
    .io_in(valid_87_io_in),
    .io_out(valid_87_io_out),
    .io_enable(valid_87_io_enable)
  );
  FF_9 valid_88 (
    .clock(valid_88_clock),
    .reset(valid_88_reset),
    .io_in(valid_88_io_in),
    .io_out(valid_88_io_out),
    .io_enable(valid_88_io_enable)
  );
  FF_9 valid_89 (
    .clock(valid_89_clock),
    .reset(valid_89_reset),
    .io_in(valid_89_io_in),
    .io_out(valid_89_io_out),
    .io_enable(valid_89_io_enable)
  );
  FF_9 valid_90 (
    .clock(valid_90_clock),
    .reset(valid_90_reset),
    .io_in(valid_90_io_in),
    .io_out(valid_90_io_out),
    .io_enable(valid_90_io_enable)
  );
  FF_9 valid_91 (
    .clock(valid_91_clock),
    .reset(valid_91_reset),
    .io_in(valid_91_io_in),
    .io_out(valid_91_io_out),
    .io_enable(valid_91_io_enable)
  );
  FF_9 valid_92 (
    .clock(valid_92_clock),
    .reset(valid_92_reset),
    .io_in(valid_92_io_in),
    .io_out(valid_92_io_out),
    .io_enable(valid_92_io_enable)
  );
  FF_9 valid_93 (
    .clock(valid_93_clock),
    .reset(valid_93_reset),
    .io_in(valid_93_io_in),
    .io_out(valid_93_io_out),
    .io_enable(valid_93_io_enable)
  );
  FF_9 valid_94 (
    .clock(valid_94_clock),
    .reset(valid_94_reset),
    .io_in(valid_94_io_in),
    .io_out(valid_94_io_out),
    .io_enable(valid_94_io_enable)
  );
  FF_9 valid_95 (
    .clock(valid_95_clock),
    .reset(valid_95_reset),
    .io_in(valid_95_io_in),
    .io_out(valid_95_io_out),
    .io_enable(valid_95_io_enable)
  );
  FF_9 valid_96 (
    .clock(valid_96_clock),
    .reset(valid_96_reset),
    .io_in(valid_96_io_in),
    .io_out(valid_96_io_out),
    .io_enable(valid_96_io_enable)
  );
  FF_9 valid_97 (
    .clock(valid_97_clock),
    .reset(valid_97_reset),
    .io_in(valid_97_io_in),
    .io_out(valid_97_io_out),
    .io_enable(valid_97_io_enable)
  );
  FF_9 valid_98 (
    .clock(valid_98_clock),
    .reset(valid_98_reset),
    .io_in(valid_98_io_in),
    .io_out(valid_98_io_out),
    .io_enable(valid_98_io_enable)
  );
  FF_9 valid_99 (
    .clock(valid_99_clock),
    .reset(valid_99_reset),
    .io_in(valid_99_io_in),
    .io_out(valid_99_io_out),
    .io_enable(valid_99_io_enable)
  );
  FF_9 valid_100 (
    .clock(valid_100_clock),
    .reset(valid_100_reset),
    .io_in(valid_100_io_in),
    .io_out(valid_100_io_out),
    .io_enable(valid_100_io_enable)
  );
  FF_9 valid_101 (
    .clock(valid_101_clock),
    .reset(valid_101_reset),
    .io_in(valid_101_io_in),
    .io_out(valid_101_io_out),
    .io_enable(valid_101_io_enable)
  );
  FF_9 valid_102 (
    .clock(valid_102_clock),
    .reset(valid_102_reset),
    .io_in(valid_102_io_in),
    .io_out(valid_102_io_out),
    .io_enable(valid_102_io_enable)
  );
  FF_9 valid_103 (
    .clock(valid_103_clock),
    .reset(valid_103_reset),
    .io_in(valid_103_io_in),
    .io_out(valid_103_io_out),
    .io_enable(valid_103_io_enable)
  );
  FF_9 valid_104 (
    .clock(valid_104_clock),
    .reset(valid_104_reset),
    .io_in(valid_104_io_in),
    .io_out(valid_104_io_out),
    .io_enable(valid_104_io_enable)
  );
  FF_9 valid_105 (
    .clock(valid_105_clock),
    .reset(valid_105_reset),
    .io_in(valid_105_io_in),
    .io_out(valid_105_io_out),
    .io_enable(valid_105_io_enable)
  );
  FF_9 valid_106 (
    .clock(valid_106_clock),
    .reset(valid_106_reset),
    .io_in(valid_106_io_in),
    .io_out(valid_106_io_out),
    .io_enable(valid_106_io_enable)
  );
  FF_9 valid_107 (
    .clock(valid_107_clock),
    .reset(valid_107_reset),
    .io_in(valid_107_io_in),
    .io_out(valid_107_io_out),
    .io_enable(valid_107_io_enable)
  );
  FF_9 valid_108 (
    .clock(valid_108_clock),
    .reset(valid_108_reset),
    .io_in(valid_108_io_in),
    .io_out(valid_108_io_out),
    .io_enable(valid_108_io_enable)
  );
  FF_9 valid_109 (
    .clock(valid_109_clock),
    .reset(valid_109_reset),
    .io_in(valid_109_io_in),
    .io_out(valid_109_io_out),
    .io_enable(valid_109_io_enable)
  );
  FF_9 valid_110 (
    .clock(valid_110_clock),
    .reset(valid_110_reset),
    .io_in(valid_110_io_in),
    .io_out(valid_110_io_out),
    .io_enable(valid_110_io_enable)
  );
  FF_9 valid_111 (
    .clock(valid_111_clock),
    .reset(valid_111_reset),
    .io_in(valid_111_io_in),
    .io_out(valid_111_io_out),
    .io_enable(valid_111_io_enable)
  );
  FF_9 valid_112 (
    .clock(valid_112_clock),
    .reset(valid_112_reset),
    .io_in(valid_112_io_in),
    .io_out(valid_112_io_out),
    .io_enable(valid_112_io_enable)
  );
  FF_9 valid_113 (
    .clock(valid_113_clock),
    .reset(valid_113_reset),
    .io_in(valid_113_io_in),
    .io_out(valid_113_io_out),
    .io_enable(valid_113_io_enable)
  );
  FF_9 valid_114 (
    .clock(valid_114_clock),
    .reset(valid_114_reset),
    .io_in(valid_114_io_in),
    .io_out(valid_114_io_out),
    .io_enable(valid_114_io_enable)
  );
  FF_9 valid_115 (
    .clock(valid_115_clock),
    .reset(valid_115_reset),
    .io_in(valid_115_io_in),
    .io_out(valid_115_io_out),
    .io_enable(valid_115_io_enable)
  );
  FF_9 valid_116 (
    .clock(valid_116_clock),
    .reset(valid_116_reset),
    .io_in(valid_116_io_in),
    .io_out(valid_116_io_out),
    .io_enable(valid_116_io_enable)
  );
  FF_9 valid_117 (
    .clock(valid_117_clock),
    .reset(valid_117_reset),
    .io_in(valid_117_io_in),
    .io_out(valid_117_io_out),
    .io_enable(valid_117_io_enable)
  );
  FF_9 valid_118 (
    .clock(valid_118_clock),
    .reset(valid_118_reset),
    .io_in(valid_118_io_in),
    .io_out(valid_118_io_out),
    .io_enable(valid_118_io_enable)
  );
  FF_9 valid_119 (
    .clock(valid_119_clock),
    .reset(valid_119_reset),
    .io_in(valid_119_io_in),
    .io_out(valid_119_io_out),
    .io_enable(valid_119_io_enable)
  );
  FF_9 valid_120 (
    .clock(valid_120_clock),
    .reset(valid_120_reset),
    .io_in(valid_120_io_in),
    .io_out(valid_120_io_out),
    .io_enable(valid_120_io_enable)
  );
  FF_9 valid_121 (
    .clock(valid_121_clock),
    .reset(valid_121_reset),
    .io_in(valid_121_io_in),
    .io_out(valid_121_io_out),
    .io_enable(valid_121_io_enable)
  );
  FF_9 valid_122 (
    .clock(valid_122_clock),
    .reset(valid_122_reset),
    .io_in(valid_122_io_in),
    .io_out(valid_122_io_out),
    .io_enable(valid_122_io_enable)
  );
  FF_9 valid_123 (
    .clock(valid_123_clock),
    .reset(valid_123_reset),
    .io_in(valid_123_io_in),
    .io_out(valid_123_io_out),
    .io_enable(valid_123_io_enable)
  );
  FF_9 valid_124 (
    .clock(valid_124_clock),
    .reset(valid_124_reset),
    .io_in(valid_124_io_in),
    .io_out(valid_124_io_out),
    .io_enable(valid_124_io_enable)
  );
  FF_9 valid_125 (
    .clock(valid_125_clock),
    .reset(valid_125_reset),
    .io_in(valid_125_io_in),
    .io_out(valid_125_io_out),
    .io_enable(valid_125_io_enable)
  );
  FF_9 valid_126 (
    .clock(valid_126_clock),
    .reset(valid_126_reset),
    .io_in(valid_126_io_in),
    .io_out(valid_126_io_out),
    .io_enable(valid_126_io_enable)
  );
  FF_9 valid_127 (
    .clock(valid_127_clock),
    .reset(valid_127_reset),
    .io_in(valid_127_io_in),
    .io_out(valid_127_io_out),
    .io_enable(valid_127_io_enable)
  );
  FF_9 valid_128 (
    .clock(valid_128_clock),
    .reset(valid_128_reset),
    .io_in(valid_128_io_in),
    .io_out(valid_128_io_out),
    .io_enable(valid_128_io_enable)
  );
  FF_9 valid_129 (
    .clock(valid_129_clock),
    .reset(valid_129_reset),
    .io_in(valid_129_io_in),
    .io_out(valid_129_io_out),
    .io_enable(valid_129_io_enable)
  );
  FF_9 valid_130 (
    .clock(valid_130_clock),
    .reset(valid_130_reset),
    .io_in(valid_130_io_in),
    .io_out(valid_130_io_out),
    .io_enable(valid_130_io_enable)
  );
  FF_9 valid_131 (
    .clock(valid_131_clock),
    .reset(valid_131_reset),
    .io_in(valid_131_io_in),
    .io_out(valid_131_io_out),
    .io_enable(valid_131_io_enable)
  );
  FF_9 valid_132 (
    .clock(valid_132_clock),
    .reset(valid_132_reset),
    .io_in(valid_132_io_in),
    .io_out(valid_132_io_out),
    .io_enable(valid_132_io_enable)
  );
  FF_9 valid_133 (
    .clock(valid_133_clock),
    .reset(valid_133_reset),
    .io_in(valid_133_io_in),
    .io_out(valid_133_io_out),
    .io_enable(valid_133_io_enable)
  );
  FF_9 valid_134 (
    .clock(valid_134_clock),
    .reset(valid_134_reset),
    .io_in(valid_134_io_in),
    .io_out(valid_134_io_out),
    .io_enable(valid_134_io_enable)
  );
  FF_9 valid_135 (
    .clock(valid_135_clock),
    .reset(valid_135_reset),
    .io_in(valid_135_io_in),
    .io_out(valid_135_io_out),
    .io_enable(valid_135_io_enable)
  );
  FF_9 valid_136 (
    .clock(valid_136_clock),
    .reset(valid_136_reset),
    .io_in(valid_136_io_in),
    .io_out(valid_136_io_out),
    .io_enable(valid_136_io_enable)
  );
  FF_9 valid_137 (
    .clock(valid_137_clock),
    .reset(valid_137_reset),
    .io_in(valid_137_io_in),
    .io_out(valid_137_io_out),
    .io_enable(valid_137_io_enable)
  );
  FF_9 valid_138 (
    .clock(valid_138_clock),
    .reset(valid_138_reset),
    .io_in(valid_138_io_in),
    .io_out(valid_138_io_out),
    .io_enable(valid_138_io_enable)
  );
  FF_9 valid_139 (
    .clock(valid_139_clock),
    .reset(valid_139_reset),
    .io_in(valid_139_io_in),
    .io_out(valid_139_io_out),
    .io_enable(valid_139_io_enable)
  );
  FF_9 valid_140 (
    .clock(valid_140_clock),
    .reset(valid_140_reset),
    .io_in(valid_140_io_in),
    .io_out(valid_140_io_out),
    .io_enable(valid_140_io_enable)
  );
  FF_9 valid_141 (
    .clock(valid_141_clock),
    .reset(valid_141_reset),
    .io_in(valid_141_io_in),
    .io_out(valid_141_io_out),
    .io_enable(valid_141_io_enable)
  );
  FF_9 valid_142 (
    .clock(valid_142_clock),
    .reset(valid_142_reset),
    .io_in(valid_142_io_in),
    .io_out(valid_142_io_out),
    .io_enable(valid_142_io_enable)
  );
  FF_9 valid_143 (
    .clock(valid_143_clock),
    .reset(valid_143_reset),
    .io_in(valid_143_io_in),
    .io_out(valid_143_io_out),
    .io_enable(valid_143_io_enable)
  );
  FF_9 valid_144 (
    .clock(valid_144_clock),
    .reset(valid_144_reset),
    .io_in(valid_144_io_in),
    .io_out(valid_144_io_out),
    .io_enable(valid_144_io_enable)
  );
  FF_9 valid_145 (
    .clock(valid_145_clock),
    .reset(valid_145_reset),
    .io_in(valid_145_io_in),
    .io_out(valid_145_io_out),
    .io_enable(valid_145_io_enable)
  );
  FF_9 valid_146 (
    .clock(valid_146_clock),
    .reset(valid_146_reset),
    .io_in(valid_146_io_in),
    .io_out(valid_146_io_out),
    .io_enable(valid_146_io_enable)
  );
  FF_9 valid_147 (
    .clock(valid_147_clock),
    .reset(valid_147_reset),
    .io_in(valid_147_io_in),
    .io_out(valid_147_io_out),
    .io_enable(valid_147_io_enable)
  );
  FF_9 valid_148 (
    .clock(valid_148_clock),
    .reset(valid_148_reset),
    .io_in(valid_148_io_in),
    .io_out(valid_148_io_out),
    .io_enable(valid_148_io_enable)
  );
  FF_9 valid_149 (
    .clock(valid_149_clock),
    .reset(valid_149_reset),
    .io_in(valid_149_io_in),
    .io_out(valid_149_io_out),
    .io_enable(valid_149_io_enable)
  );
  FF_9 valid_150 (
    .clock(valid_150_clock),
    .reset(valid_150_reset),
    .io_in(valid_150_io_in),
    .io_out(valid_150_io_out),
    .io_enable(valid_150_io_enable)
  );
  FF_9 valid_151 (
    .clock(valid_151_clock),
    .reset(valid_151_reset),
    .io_in(valid_151_io_in),
    .io_out(valid_151_io_out),
    .io_enable(valid_151_io_enable)
  );
  FF_9 valid_152 (
    .clock(valid_152_clock),
    .reset(valid_152_reset),
    .io_in(valid_152_io_in),
    .io_out(valid_152_io_out),
    .io_enable(valid_152_io_enable)
  );
  FF_9 valid_153 (
    .clock(valid_153_clock),
    .reset(valid_153_reset),
    .io_in(valid_153_io_in),
    .io_out(valid_153_io_out),
    .io_enable(valid_153_io_enable)
  );
  FF_9 valid_154 (
    .clock(valid_154_clock),
    .reset(valid_154_reset),
    .io_in(valid_154_io_in),
    .io_out(valid_154_io_out),
    .io_enable(valid_154_io_enable)
  );
  FF_9 valid_155 (
    .clock(valid_155_clock),
    .reset(valid_155_reset),
    .io_in(valid_155_io_in),
    .io_out(valid_155_io_out),
    .io_enable(valid_155_io_enable)
  );
  FF_9 valid_156 (
    .clock(valid_156_clock),
    .reset(valid_156_reset),
    .io_in(valid_156_io_in),
    .io_out(valid_156_io_out),
    .io_enable(valid_156_io_enable)
  );
  FF_9 valid_157 (
    .clock(valid_157_clock),
    .reset(valid_157_reset),
    .io_in(valid_157_io_in),
    .io_out(valid_157_io_out),
    .io_enable(valid_157_io_enable)
  );
  FF_9 valid_158 (
    .clock(valid_158_clock),
    .reset(valid_158_reset),
    .io_in(valid_158_io_in),
    .io_out(valid_158_io_out),
    .io_enable(valid_158_io_enable)
  );
  FF_9 valid_159 (
    .clock(valid_159_clock),
    .reset(valid_159_reset),
    .io_in(valid_159_io_in),
    .io_out(valid_159_io_out),
    .io_enable(valid_159_io_enable)
  );
  FF_9 valid_160 (
    .clock(valid_160_clock),
    .reset(valid_160_reset),
    .io_in(valid_160_io_in),
    .io_out(valid_160_io_out),
    .io_enable(valid_160_io_enable)
  );
  FF_9 valid_161 (
    .clock(valid_161_clock),
    .reset(valid_161_reset),
    .io_in(valid_161_io_in),
    .io_out(valid_161_io_out),
    .io_enable(valid_161_io_enable)
  );
  FF_9 valid_162 (
    .clock(valid_162_clock),
    .reset(valid_162_reset),
    .io_in(valid_162_io_in),
    .io_out(valid_162_io_out),
    .io_enable(valid_162_io_enable)
  );
  FF_9 valid_163 (
    .clock(valid_163_clock),
    .reset(valid_163_reset),
    .io_in(valid_163_io_in),
    .io_out(valid_163_io_out),
    .io_enable(valid_163_io_enable)
  );
  FF_9 valid_164 (
    .clock(valid_164_clock),
    .reset(valid_164_reset),
    .io_in(valid_164_io_in),
    .io_out(valid_164_io_out),
    .io_enable(valid_164_io_enable)
  );
  FF_9 valid_165 (
    .clock(valid_165_clock),
    .reset(valid_165_reset),
    .io_in(valid_165_io_in),
    .io_out(valid_165_io_out),
    .io_enable(valid_165_io_enable)
  );
  FF_9 valid_166 (
    .clock(valid_166_clock),
    .reset(valid_166_reset),
    .io_in(valid_166_io_in),
    .io_out(valid_166_io_out),
    .io_enable(valid_166_io_enable)
  );
  FF_9 valid_167 (
    .clock(valid_167_clock),
    .reset(valid_167_reset),
    .io_in(valid_167_io_in),
    .io_out(valid_167_io_out),
    .io_enable(valid_167_io_enable)
  );
  FF_9 valid_168 (
    .clock(valid_168_clock),
    .reset(valid_168_reset),
    .io_in(valid_168_io_in),
    .io_out(valid_168_io_out),
    .io_enable(valid_168_io_enable)
  );
  FF_9 valid_169 (
    .clock(valid_169_clock),
    .reset(valid_169_reset),
    .io_in(valid_169_io_in),
    .io_out(valid_169_io_out),
    .io_enable(valid_169_io_enable)
  );
  FF_9 valid_170 (
    .clock(valid_170_clock),
    .reset(valid_170_reset),
    .io_in(valid_170_io_in),
    .io_out(valid_170_io_out),
    .io_enable(valid_170_io_enable)
  );
  FF_9 valid_171 (
    .clock(valid_171_clock),
    .reset(valid_171_reset),
    .io_in(valid_171_io_in),
    .io_out(valid_171_io_out),
    .io_enable(valid_171_io_enable)
  );
  FF_9 valid_172 (
    .clock(valid_172_clock),
    .reset(valid_172_reset),
    .io_in(valid_172_io_in),
    .io_out(valid_172_io_out),
    .io_enable(valid_172_io_enable)
  );
  FF_9 valid_173 (
    .clock(valid_173_clock),
    .reset(valid_173_reset),
    .io_in(valid_173_io_in),
    .io_out(valid_173_io_out),
    .io_enable(valid_173_io_enable)
  );
  FF_9 valid_174 (
    .clock(valid_174_clock),
    .reset(valid_174_reset),
    .io_in(valid_174_io_in),
    .io_out(valid_174_io_out),
    .io_enable(valid_174_io_enable)
  );
  FF_9 valid_175 (
    .clock(valid_175_clock),
    .reset(valid_175_reset),
    .io_in(valid_175_io_in),
    .io_out(valid_175_io_out),
    .io_enable(valid_175_io_enable)
  );
  FF_9 valid_176 (
    .clock(valid_176_clock),
    .reset(valid_176_reset),
    .io_in(valid_176_io_in),
    .io_out(valid_176_io_out),
    .io_enable(valid_176_io_enable)
  );
  FF_9 valid_177 (
    .clock(valid_177_clock),
    .reset(valid_177_reset),
    .io_in(valid_177_io_in),
    .io_out(valid_177_io_out),
    .io_enable(valid_177_io_enable)
  );
  FF_9 valid_178 (
    .clock(valid_178_clock),
    .reset(valid_178_reset),
    .io_in(valid_178_io_in),
    .io_out(valid_178_io_out),
    .io_enable(valid_178_io_enable)
  );
  FF_9 valid_179 (
    .clock(valid_179_clock),
    .reset(valid_179_reset),
    .io_in(valid_179_io_in),
    .io_out(valid_179_io_out),
    .io_enable(valid_179_io_enable)
  );
  FF_9 valid_180 (
    .clock(valid_180_clock),
    .reset(valid_180_reset),
    .io_in(valid_180_io_in),
    .io_out(valid_180_io_out),
    .io_enable(valid_180_io_enable)
  );
  FF_9 valid_181 (
    .clock(valid_181_clock),
    .reset(valid_181_reset),
    .io_in(valid_181_io_in),
    .io_out(valid_181_io_out),
    .io_enable(valid_181_io_enable)
  );
  FF_9 valid_182 (
    .clock(valid_182_clock),
    .reset(valid_182_reset),
    .io_in(valid_182_io_in),
    .io_out(valid_182_io_out),
    .io_enable(valid_182_io_enable)
  );
  FF_9 valid_183 (
    .clock(valid_183_clock),
    .reset(valid_183_reset),
    .io_in(valid_183_io_in),
    .io_out(valid_183_io_out),
    .io_enable(valid_183_io_enable)
  );
  FF_9 valid_184 (
    .clock(valid_184_clock),
    .reset(valid_184_reset),
    .io_in(valid_184_io_in),
    .io_out(valid_184_io_out),
    .io_enable(valid_184_io_enable)
  );
  FF_9 valid_185 (
    .clock(valid_185_clock),
    .reset(valid_185_reset),
    .io_in(valid_185_io_in),
    .io_out(valid_185_io_out),
    .io_enable(valid_185_io_enable)
  );
  FF_9 valid_186 (
    .clock(valid_186_clock),
    .reset(valid_186_reset),
    .io_in(valid_186_io_in),
    .io_out(valid_186_io_out),
    .io_enable(valid_186_io_enable)
  );
  FF_9 valid_187 (
    .clock(valid_187_clock),
    .reset(valid_187_reset),
    .io_in(valid_187_io_in),
    .io_out(valid_187_io_out),
    .io_enable(valid_187_io_enable)
  );
  FF_9 valid_188 (
    .clock(valid_188_clock),
    .reset(valid_188_reset),
    .io_in(valid_188_io_in),
    .io_out(valid_188_io_out),
    .io_enable(valid_188_io_enable)
  );
  FF_9 valid_189 (
    .clock(valid_189_clock),
    .reset(valid_189_reset),
    .io_in(valid_189_io_in),
    .io_out(valid_189_io_out),
    .io_enable(valid_189_io_enable)
  );
  FF_9 valid_190 (
    .clock(valid_190_clock),
    .reset(valid_190_reset),
    .io_in(valid_190_io_in),
    .io_out(valid_190_io_out),
    .io_enable(valid_190_io_enable)
  );
  FF_9 valid_191 (
    .clock(valid_191_clock),
    .reset(valid_191_reset),
    .io_in(valid_191_io_in),
    .io_out(valid_191_io_out),
    .io_enable(valid_191_io_enable)
  );
  FF_9 valid_192 (
    .clock(valid_192_clock),
    .reset(valid_192_reset),
    .io_in(valid_192_io_in),
    .io_out(valid_192_io_out),
    .io_enable(valid_192_io_enable)
  );
  FF_9 valid_193 (
    .clock(valid_193_clock),
    .reset(valid_193_reset),
    .io_in(valid_193_io_in),
    .io_out(valid_193_io_out),
    .io_enable(valid_193_io_enable)
  );
  FF_9 valid_194 (
    .clock(valid_194_clock),
    .reset(valid_194_reset),
    .io_in(valid_194_io_in),
    .io_out(valid_194_io_out),
    .io_enable(valid_194_io_enable)
  );
  FF_9 valid_195 (
    .clock(valid_195_clock),
    .reset(valid_195_reset),
    .io_in(valid_195_io_in),
    .io_out(valid_195_io_out),
    .io_enable(valid_195_io_enable)
  );
  FF_9 valid_196 (
    .clock(valid_196_clock),
    .reset(valid_196_reset),
    .io_in(valid_196_io_in),
    .io_out(valid_196_io_out),
    .io_enable(valid_196_io_enable)
  );
  FF_9 valid_197 (
    .clock(valid_197_clock),
    .reset(valid_197_reset),
    .io_in(valid_197_io_in),
    .io_out(valid_197_io_out),
    .io_enable(valid_197_io_enable)
  );
  FF_9 valid_198 (
    .clock(valid_198_clock),
    .reset(valid_198_reset),
    .io_in(valid_198_io_in),
    .io_out(valid_198_io_out),
    .io_enable(valid_198_io_enable)
  );
  FF_9 valid_199 (
    .clock(valid_199_clock),
    .reset(valid_199_reset),
    .io_in(valid_199_io_in),
    .io_out(valid_199_io_out),
    .io_enable(valid_199_io_enable)
  );
  FF_9 valid_200 (
    .clock(valid_200_clock),
    .reset(valid_200_reset),
    .io_in(valid_200_io_in),
    .io_out(valid_200_io_out),
    .io_enable(valid_200_io_enable)
  );
  FF_9 valid_201 (
    .clock(valid_201_clock),
    .reset(valid_201_reset),
    .io_in(valid_201_io_in),
    .io_out(valid_201_io_out),
    .io_enable(valid_201_io_enable)
  );
  FF_9 valid_202 (
    .clock(valid_202_clock),
    .reset(valid_202_reset),
    .io_in(valid_202_io_in),
    .io_out(valid_202_io_out),
    .io_enable(valid_202_io_enable)
  );
  FF_9 valid_203 (
    .clock(valid_203_clock),
    .reset(valid_203_reset),
    .io_in(valid_203_io_in),
    .io_out(valid_203_io_out),
    .io_enable(valid_203_io_enable)
  );
  FF_9 valid_204 (
    .clock(valid_204_clock),
    .reset(valid_204_reset),
    .io_in(valid_204_io_in),
    .io_out(valid_204_io_out),
    .io_enable(valid_204_io_enable)
  );
  FF_9 valid_205 (
    .clock(valid_205_clock),
    .reset(valid_205_reset),
    .io_in(valid_205_io_in),
    .io_out(valid_205_io_out),
    .io_enable(valid_205_io_enable)
  );
  FF_9 valid_206 (
    .clock(valid_206_clock),
    .reset(valid_206_reset),
    .io_in(valid_206_io_in),
    .io_out(valid_206_io_out),
    .io_enable(valid_206_io_enable)
  );
  FF_9 valid_207 (
    .clock(valid_207_clock),
    .reset(valid_207_reset),
    .io_in(valid_207_io_in),
    .io_out(valid_207_io_out),
    .io_enable(valid_207_io_enable)
  );
  FF_9 valid_208 (
    .clock(valid_208_clock),
    .reset(valid_208_reset),
    .io_in(valid_208_io_in),
    .io_out(valid_208_io_out),
    .io_enable(valid_208_io_enable)
  );
  FF_9 valid_209 (
    .clock(valid_209_clock),
    .reset(valid_209_reset),
    .io_in(valid_209_io_in),
    .io_out(valid_209_io_out),
    .io_enable(valid_209_io_enable)
  );
  FF_9 valid_210 (
    .clock(valid_210_clock),
    .reset(valid_210_reset),
    .io_in(valid_210_io_in),
    .io_out(valid_210_io_out),
    .io_enable(valid_210_io_enable)
  );
  FF_9 valid_211 (
    .clock(valid_211_clock),
    .reset(valid_211_reset),
    .io_in(valid_211_io_in),
    .io_out(valid_211_io_out),
    .io_enable(valid_211_io_enable)
  );
  FF_9 valid_212 (
    .clock(valid_212_clock),
    .reset(valid_212_reset),
    .io_in(valid_212_io_in),
    .io_out(valid_212_io_out),
    .io_enable(valid_212_io_enable)
  );
  FF_9 valid_213 (
    .clock(valid_213_clock),
    .reset(valid_213_reset),
    .io_in(valid_213_io_in),
    .io_out(valid_213_io_out),
    .io_enable(valid_213_io_enable)
  );
  FF_9 valid_214 (
    .clock(valid_214_clock),
    .reset(valid_214_reset),
    .io_in(valid_214_io_in),
    .io_out(valid_214_io_out),
    .io_enable(valid_214_io_enable)
  );
  FF_9 valid_215 (
    .clock(valid_215_clock),
    .reset(valid_215_reset),
    .io_in(valid_215_io_in),
    .io_out(valid_215_io_out),
    .io_enable(valid_215_io_enable)
  );
  FF_9 valid_216 (
    .clock(valid_216_clock),
    .reset(valid_216_reset),
    .io_in(valid_216_io_in),
    .io_out(valid_216_io_out),
    .io_enable(valid_216_io_enable)
  );
  FF_9 valid_217 (
    .clock(valid_217_clock),
    .reset(valid_217_reset),
    .io_in(valid_217_io_in),
    .io_out(valid_217_io_out),
    .io_enable(valid_217_io_enable)
  );
  FF_9 valid_218 (
    .clock(valid_218_clock),
    .reset(valid_218_reset),
    .io_in(valid_218_io_in),
    .io_out(valid_218_io_out),
    .io_enable(valid_218_io_enable)
  );
  FF_9 valid_219 (
    .clock(valid_219_clock),
    .reset(valid_219_reset),
    .io_in(valid_219_io_in),
    .io_out(valid_219_io_out),
    .io_enable(valid_219_io_enable)
  );
  FF_9 valid_220 (
    .clock(valid_220_clock),
    .reset(valid_220_reset),
    .io_in(valid_220_io_in),
    .io_out(valid_220_io_out),
    .io_enable(valid_220_io_enable)
  );
  FF_9 valid_221 (
    .clock(valid_221_clock),
    .reset(valid_221_reset),
    .io_in(valid_221_io_in),
    .io_out(valid_221_io_out),
    .io_enable(valid_221_io_enable)
  );
  FF_9 valid_222 (
    .clock(valid_222_clock),
    .reset(valid_222_reset),
    .io_in(valid_222_io_in),
    .io_out(valid_222_io_out),
    .io_enable(valid_222_io_enable)
  );
  FF_9 valid_223 (
    .clock(valid_223_clock),
    .reset(valid_223_reset),
    .io_in(valid_223_io_in),
    .io_out(valid_223_io_out),
    .io_enable(valid_223_io_enable)
  );
  FF_9 valid_224 (
    .clock(valid_224_clock),
    .reset(valid_224_reset),
    .io_in(valid_224_io_in),
    .io_out(valid_224_io_out),
    .io_enable(valid_224_io_enable)
  );
  FF_9 valid_225 (
    .clock(valid_225_clock),
    .reset(valid_225_reset),
    .io_in(valid_225_io_in),
    .io_out(valid_225_io_out),
    .io_enable(valid_225_io_enable)
  );
  FF_9 valid_226 (
    .clock(valid_226_clock),
    .reset(valid_226_reset),
    .io_in(valid_226_io_in),
    .io_out(valid_226_io_out),
    .io_enable(valid_226_io_enable)
  );
  FF_9 valid_227 (
    .clock(valid_227_clock),
    .reset(valid_227_reset),
    .io_in(valid_227_io_in),
    .io_out(valid_227_io_out),
    .io_enable(valid_227_io_enable)
  );
  FF_9 valid_228 (
    .clock(valid_228_clock),
    .reset(valid_228_reset),
    .io_in(valid_228_io_in),
    .io_out(valid_228_io_out),
    .io_enable(valid_228_io_enable)
  );
  FF_9 valid_229 (
    .clock(valid_229_clock),
    .reset(valid_229_reset),
    .io_in(valid_229_io_in),
    .io_out(valid_229_io_out),
    .io_enable(valid_229_io_enable)
  );
  FF_9 valid_230 (
    .clock(valid_230_clock),
    .reset(valid_230_reset),
    .io_in(valid_230_io_in),
    .io_out(valid_230_io_out),
    .io_enable(valid_230_io_enable)
  );
  FF_9 valid_231 (
    .clock(valid_231_clock),
    .reset(valid_231_reset),
    .io_in(valid_231_io_in),
    .io_out(valid_231_io_out),
    .io_enable(valid_231_io_enable)
  );
  FF_9 valid_232 (
    .clock(valid_232_clock),
    .reset(valid_232_reset),
    .io_in(valid_232_io_in),
    .io_out(valid_232_io_out),
    .io_enable(valid_232_io_enable)
  );
  FF_9 valid_233 (
    .clock(valid_233_clock),
    .reset(valid_233_reset),
    .io_in(valid_233_io_in),
    .io_out(valid_233_io_out),
    .io_enable(valid_233_io_enable)
  );
  FF_9 valid_234 (
    .clock(valid_234_clock),
    .reset(valid_234_reset),
    .io_in(valid_234_io_in),
    .io_out(valid_234_io_out),
    .io_enable(valid_234_io_enable)
  );
  FF_9 valid_235 (
    .clock(valid_235_clock),
    .reset(valid_235_reset),
    .io_in(valid_235_io_in),
    .io_out(valid_235_io_out),
    .io_enable(valid_235_io_enable)
  );
  FF_9 valid_236 (
    .clock(valid_236_clock),
    .reset(valid_236_reset),
    .io_in(valid_236_io_in),
    .io_out(valid_236_io_out),
    .io_enable(valid_236_io_enable)
  );
  FF_9 valid_237 (
    .clock(valid_237_clock),
    .reset(valid_237_reset),
    .io_in(valid_237_io_in),
    .io_out(valid_237_io_out),
    .io_enable(valid_237_io_enable)
  );
  FF_9 valid_238 (
    .clock(valid_238_clock),
    .reset(valid_238_reset),
    .io_in(valid_238_io_in),
    .io_out(valid_238_io_out),
    .io_enable(valid_238_io_enable)
  );
  FF_9 valid_239 (
    .clock(valid_239_clock),
    .reset(valid_239_reset),
    .io_in(valid_239_io_in),
    .io_out(valid_239_io_out),
    .io_enable(valid_239_io_enable)
  );
  FF_9 valid_240 (
    .clock(valid_240_clock),
    .reset(valid_240_reset),
    .io_in(valid_240_io_in),
    .io_out(valid_240_io_out),
    .io_enable(valid_240_io_enable)
  );
  FF_9 valid_241 (
    .clock(valid_241_clock),
    .reset(valid_241_reset),
    .io_in(valid_241_io_in),
    .io_out(valid_241_io_out),
    .io_enable(valid_241_io_enable)
  );
  FF_9 valid_242 (
    .clock(valid_242_clock),
    .reset(valid_242_reset),
    .io_in(valid_242_io_in),
    .io_out(valid_242_io_out),
    .io_enable(valid_242_io_enable)
  );
  FF_9 valid_243 (
    .clock(valid_243_clock),
    .reset(valid_243_reset),
    .io_in(valid_243_io_in),
    .io_out(valid_243_io_out),
    .io_enable(valid_243_io_enable)
  );
  FF_9 valid_244 (
    .clock(valid_244_clock),
    .reset(valid_244_reset),
    .io_in(valid_244_io_in),
    .io_out(valid_244_io_out),
    .io_enable(valid_244_io_enable)
  );
  FF_9 valid_245 (
    .clock(valid_245_clock),
    .reset(valid_245_reset),
    .io_in(valid_245_io_in),
    .io_out(valid_245_io_out),
    .io_enable(valid_245_io_enable)
  );
  FF_9 valid_246 (
    .clock(valid_246_clock),
    .reset(valid_246_reset),
    .io_in(valid_246_io_in),
    .io_out(valid_246_io_out),
    .io_enable(valid_246_io_enable)
  );
  FF_9 valid_247 (
    .clock(valid_247_clock),
    .reset(valid_247_reset),
    .io_in(valid_247_io_in),
    .io_out(valid_247_io_out),
    .io_enable(valid_247_io_enable)
  );
  FF_9 valid_248 (
    .clock(valid_248_clock),
    .reset(valid_248_reset),
    .io_in(valid_248_io_in),
    .io_out(valid_248_io_out),
    .io_enable(valid_248_io_enable)
  );
  FF_9 valid_249 (
    .clock(valid_249_clock),
    .reset(valid_249_reset),
    .io_in(valid_249_io_in),
    .io_out(valid_249_io_out),
    .io_enable(valid_249_io_enable)
  );
  FF_9 valid_250 (
    .clock(valid_250_clock),
    .reset(valid_250_reset),
    .io_in(valid_250_io_in),
    .io_out(valid_250_io_out),
    .io_enable(valid_250_io_enable)
  );
  FF_9 valid_251 (
    .clock(valid_251_clock),
    .reset(valid_251_reset),
    .io_in(valid_251_io_in),
    .io_out(valid_251_io_out),
    .io_enable(valid_251_io_enable)
  );
  FF_9 valid_252 (
    .clock(valid_252_clock),
    .reset(valid_252_reset),
    .io_in(valid_252_io_in),
    .io_out(valid_252_io_out),
    .io_enable(valid_252_io_enable)
  );
  FF_9 valid_253 (
    .clock(valid_253_clock),
    .reset(valid_253_reset),
    .io_in(valid_253_io_in),
    .io_out(valid_253_io_out),
    .io_enable(valid_253_io_enable)
  );
  FF_9 valid_254 (
    .clock(valid_254_clock),
    .reset(valid_254_reset),
    .io_in(valid_254_io_in),
    .io_out(valid_254_io_out),
    .io_enable(valid_254_io_enable)
  );
  FF_9 valid_255 (
    .clock(valid_255_clock),
    .reset(valid_255_reset),
    .io_in(valid_255_io_in),
    .io_out(valid_255_io_out),
    .io_enable(valid_255_io_enable)
  );
  FF_9 valid_256 (
    .clock(valid_256_clock),
    .reset(valid_256_reset),
    .io_in(valid_256_io_in),
    .io_out(valid_256_io_out),
    .io_enable(valid_256_io_enable)
  );
  FF_9 valid_257 (
    .clock(valid_257_clock),
    .reset(valid_257_reset),
    .io_in(valid_257_io_in),
    .io_out(valid_257_io_out),
    .io_enable(valid_257_io_enable)
  );
  FF_9 valid_258 (
    .clock(valid_258_clock),
    .reset(valid_258_reset),
    .io_in(valid_258_io_in),
    .io_out(valid_258_io_out),
    .io_enable(valid_258_io_enable)
  );
  FF_9 valid_259 (
    .clock(valid_259_clock),
    .reset(valid_259_reset),
    .io_in(valid_259_io_in),
    .io_out(valid_259_io_out),
    .io_enable(valid_259_io_enable)
  );
  FF_9 valid_260 (
    .clock(valid_260_clock),
    .reset(valid_260_reset),
    .io_in(valid_260_io_in),
    .io_out(valid_260_io_out),
    .io_enable(valid_260_io_enable)
  );
  FF_9 valid_261 (
    .clock(valid_261_clock),
    .reset(valid_261_reset),
    .io_in(valid_261_io_in),
    .io_out(valid_261_io_out),
    .io_enable(valid_261_io_enable)
  );
  FF_9 valid_262 (
    .clock(valid_262_clock),
    .reset(valid_262_reset),
    .io_in(valid_262_io_in),
    .io_out(valid_262_io_out),
    .io_enable(valid_262_io_enable)
  );
  FF_9 valid_263 (
    .clock(valid_263_clock),
    .reset(valid_263_reset),
    .io_in(valid_263_io_in),
    .io_out(valid_263_io_out),
    .io_enable(valid_263_io_enable)
  );
  FF_9 valid_264 (
    .clock(valid_264_clock),
    .reset(valid_264_reset),
    .io_in(valid_264_io_in),
    .io_out(valid_264_io_out),
    .io_enable(valid_264_io_enable)
  );
  FF_9 valid_265 (
    .clock(valid_265_clock),
    .reset(valid_265_reset),
    .io_in(valid_265_io_in),
    .io_out(valid_265_io_out),
    .io_enable(valid_265_io_enable)
  );
  FF_9 valid_266 (
    .clock(valid_266_clock),
    .reset(valid_266_reset),
    .io_in(valid_266_io_in),
    .io_out(valid_266_io_out),
    .io_enable(valid_266_io_enable)
  );
  FF_9 valid_267 (
    .clock(valid_267_clock),
    .reset(valid_267_reset),
    .io_in(valid_267_io_in),
    .io_out(valid_267_io_out),
    .io_enable(valid_267_io_enable)
  );
  FF_9 valid_268 (
    .clock(valid_268_clock),
    .reset(valid_268_reset),
    .io_in(valid_268_io_in),
    .io_out(valid_268_io_out),
    .io_enable(valid_268_io_enable)
  );
  FF_9 valid_269 (
    .clock(valid_269_clock),
    .reset(valid_269_reset),
    .io_in(valid_269_io_in),
    .io_out(valid_269_io_out),
    .io_enable(valid_269_io_enable)
  );
  FF_9 valid_270 (
    .clock(valid_270_clock),
    .reset(valid_270_reset),
    .io_in(valid_270_io_in),
    .io_out(valid_270_io_out),
    .io_enable(valid_270_io_enable)
  );
  FF_9 valid_271 (
    .clock(valid_271_clock),
    .reset(valid_271_reset),
    .io_in(valid_271_io_in),
    .io_out(valid_271_io_out),
    .io_enable(valid_271_io_enable)
  );
  FF_9 valid_272 (
    .clock(valid_272_clock),
    .reset(valid_272_reset),
    .io_in(valid_272_io_in),
    .io_out(valid_272_io_out),
    .io_enable(valid_272_io_enable)
  );
  FF_9 valid_273 (
    .clock(valid_273_clock),
    .reset(valid_273_reset),
    .io_in(valid_273_io_in),
    .io_out(valid_273_io_out),
    .io_enable(valid_273_io_enable)
  );
  FF_9 valid_274 (
    .clock(valid_274_clock),
    .reset(valid_274_reset),
    .io_in(valid_274_io_in),
    .io_out(valid_274_io_out),
    .io_enable(valid_274_io_enable)
  );
  FF_9 valid_275 (
    .clock(valid_275_clock),
    .reset(valid_275_reset),
    .io_in(valid_275_io_in),
    .io_out(valid_275_io_out),
    .io_enable(valid_275_io_enable)
  );
  FF_9 valid_276 (
    .clock(valid_276_clock),
    .reset(valid_276_reset),
    .io_in(valid_276_io_in),
    .io_out(valid_276_io_out),
    .io_enable(valid_276_io_enable)
  );
  FF_9 valid_277 (
    .clock(valid_277_clock),
    .reset(valid_277_reset),
    .io_in(valid_277_io_in),
    .io_out(valid_277_io_out),
    .io_enable(valid_277_io_enable)
  );
  FF_9 valid_278 (
    .clock(valid_278_clock),
    .reset(valid_278_reset),
    .io_in(valid_278_io_in),
    .io_out(valid_278_io_out),
    .io_enable(valid_278_io_enable)
  );
  FF_9 valid_279 (
    .clock(valid_279_clock),
    .reset(valid_279_reset),
    .io_in(valid_279_io_in),
    .io_out(valid_279_io_out),
    .io_enable(valid_279_io_enable)
  );
  FF_9 valid_280 (
    .clock(valid_280_clock),
    .reset(valid_280_reset),
    .io_in(valid_280_io_in),
    .io_out(valid_280_io_out),
    .io_enable(valid_280_io_enable)
  );
  FF_9 valid_281 (
    .clock(valid_281_clock),
    .reset(valid_281_reset),
    .io_in(valid_281_io_in),
    .io_out(valid_281_io_out),
    .io_enable(valid_281_io_enable)
  );
  FF_9 valid_282 (
    .clock(valid_282_clock),
    .reset(valid_282_reset),
    .io_in(valid_282_io_in),
    .io_out(valid_282_io_out),
    .io_enable(valid_282_io_enable)
  );
  FF_9 valid_283 (
    .clock(valid_283_clock),
    .reset(valid_283_reset),
    .io_in(valid_283_io_in),
    .io_out(valid_283_io_out),
    .io_enable(valid_283_io_enable)
  );
  FF_9 valid_284 (
    .clock(valid_284_clock),
    .reset(valid_284_reset),
    .io_in(valid_284_io_in),
    .io_out(valid_284_io_out),
    .io_enable(valid_284_io_enable)
  );
  FF_9 valid_285 (
    .clock(valid_285_clock),
    .reset(valid_285_reset),
    .io_in(valid_285_io_in),
    .io_out(valid_285_io_out),
    .io_enable(valid_285_io_enable)
  );
  FF_9 valid_286 (
    .clock(valid_286_clock),
    .reset(valid_286_reset),
    .io_in(valid_286_io_in),
    .io_out(valid_286_io_out),
    .io_enable(valid_286_io_enable)
  );
  FF_9 valid_287 (
    .clock(valid_287_clock),
    .reset(valid_287_reset),
    .io_in(valid_287_io_in),
    .io_out(valid_287_io_out),
    .io_enable(valid_287_io_enable)
  );
  FF_9 valid_288 (
    .clock(valid_288_clock),
    .reset(valid_288_reset),
    .io_in(valid_288_io_in),
    .io_out(valid_288_io_out),
    .io_enable(valid_288_io_enable)
  );
  FF_9 valid_289 (
    .clock(valid_289_clock),
    .reset(valid_289_reset),
    .io_in(valid_289_io_in),
    .io_out(valid_289_io_out),
    .io_enable(valid_289_io_enable)
  );
  FF_9 valid_290 (
    .clock(valid_290_clock),
    .reset(valid_290_reset),
    .io_in(valid_290_io_in),
    .io_out(valid_290_io_out),
    .io_enable(valid_290_io_enable)
  );
  FF_9 valid_291 (
    .clock(valid_291_clock),
    .reset(valid_291_reset),
    .io_in(valid_291_io_in),
    .io_out(valid_291_io_out),
    .io_enable(valid_291_io_enable)
  );
  FF_9 valid_292 (
    .clock(valid_292_clock),
    .reset(valid_292_reset),
    .io_in(valid_292_io_in),
    .io_out(valid_292_io_out),
    .io_enable(valid_292_io_enable)
  );
  FF_9 valid_293 (
    .clock(valid_293_clock),
    .reset(valid_293_reset),
    .io_in(valid_293_io_in),
    .io_out(valid_293_io_out),
    .io_enable(valid_293_io_enable)
  );
  FF_9 valid_294 (
    .clock(valid_294_clock),
    .reset(valid_294_reset),
    .io_in(valid_294_io_in),
    .io_out(valid_294_io_out),
    .io_enable(valid_294_io_enable)
  );
  FF_9 valid_295 (
    .clock(valid_295_clock),
    .reset(valid_295_reset),
    .io_in(valid_295_io_in),
    .io_out(valid_295_io_out),
    .io_enable(valid_295_io_enable)
  );
  FF_9 valid_296 (
    .clock(valid_296_clock),
    .reset(valid_296_reset),
    .io_in(valid_296_io_in),
    .io_out(valid_296_io_out),
    .io_enable(valid_296_io_enable)
  );
  FF_9 valid_297 (
    .clock(valid_297_clock),
    .reset(valid_297_reset),
    .io_in(valid_297_io_in),
    .io_out(valid_297_io_out),
    .io_enable(valid_297_io_enable)
  );
  FF_9 valid_298 (
    .clock(valid_298_clock),
    .reset(valid_298_reset),
    .io_in(valid_298_io_in),
    .io_out(valid_298_io_out),
    .io_enable(valid_298_io_enable)
  );
  FF_9 valid_299 (
    .clock(valid_299_clock),
    .reset(valid_299_reset),
    .io_in(valid_299_io_in),
    .io_out(valid_299_io_out),
    .io_enable(valid_299_io_enable)
  );
  FF_9 valid_300 (
    .clock(valid_300_clock),
    .reset(valid_300_reset),
    .io_in(valid_300_io_in),
    .io_out(valid_300_io_out),
    .io_enable(valid_300_io_enable)
  );
  FF_9 valid_301 (
    .clock(valid_301_clock),
    .reset(valid_301_reset),
    .io_in(valid_301_io_in),
    .io_out(valid_301_io_out),
    .io_enable(valid_301_io_enable)
  );
  FF_9 valid_302 (
    .clock(valid_302_clock),
    .reset(valid_302_reset),
    .io_in(valid_302_io_in),
    .io_out(valid_302_io_out),
    .io_enable(valid_302_io_enable)
  );
  FF_9 valid_303 (
    .clock(valid_303_clock),
    .reset(valid_303_reset),
    .io_in(valid_303_io_in),
    .io_out(valid_303_io_out),
    .io_enable(valid_303_io_enable)
  );
  FF_9 valid_304 (
    .clock(valid_304_clock),
    .reset(valid_304_reset),
    .io_in(valid_304_io_in),
    .io_out(valid_304_io_out),
    .io_enable(valid_304_io_enable)
  );
  FF_9 valid_305 (
    .clock(valid_305_clock),
    .reset(valid_305_reset),
    .io_in(valid_305_io_in),
    .io_out(valid_305_io_out),
    .io_enable(valid_305_io_enable)
  );
  FF_9 valid_306 (
    .clock(valid_306_clock),
    .reset(valid_306_reset),
    .io_in(valid_306_io_in),
    .io_out(valid_306_io_out),
    .io_enable(valid_306_io_enable)
  );
  FF_9 valid_307 (
    .clock(valid_307_clock),
    .reset(valid_307_reset),
    .io_in(valid_307_io_in),
    .io_out(valid_307_io_out),
    .io_enable(valid_307_io_enable)
  );
  FF_9 valid_308 (
    .clock(valid_308_clock),
    .reset(valid_308_reset),
    .io_in(valid_308_io_in),
    .io_out(valid_308_io_out),
    .io_enable(valid_308_io_enable)
  );
  FF_9 valid_309 (
    .clock(valid_309_clock),
    .reset(valid_309_reset),
    .io_in(valid_309_io_in),
    .io_out(valid_309_io_out),
    .io_enable(valid_309_io_enable)
  );
  FF_9 valid_310 (
    .clock(valid_310_clock),
    .reset(valid_310_reset),
    .io_in(valid_310_io_in),
    .io_out(valid_310_io_out),
    .io_enable(valid_310_io_enable)
  );
  FF_9 valid_311 (
    .clock(valid_311_clock),
    .reset(valid_311_reset),
    .io_in(valid_311_io_in),
    .io_out(valid_311_io_out),
    .io_enable(valid_311_io_enable)
  );
  FF_9 valid_312 (
    .clock(valid_312_clock),
    .reset(valid_312_reset),
    .io_in(valid_312_io_in),
    .io_out(valid_312_io_out),
    .io_enable(valid_312_io_enable)
  );
  FF_9 valid_313 (
    .clock(valid_313_clock),
    .reset(valid_313_reset),
    .io_in(valid_313_io_in),
    .io_out(valid_313_io_out),
    .io_enable(valid_313_io_enable)
  );
  FF_9 valid_314 (
    .clock(valid_314_clock),
    .reset(valid_314_reset),
    .io_in(valid_314_io_in),
    .io_out(valid_314_io_out),
    .io_enable(valid_314_io_enable)
  );
  FF_9 valid_315 (
    .clock(valid_315_clock),
    .reset(valid_315_reset),
    .io_in(valid_315_io_in),
    .io_out(valid_315_io_out),
    .io_enable(valid_315_io_enable)
  );
  FF_9 valid_316 (
    .clock(valid_316_clock),
    .reset(valid_316_reset),
    .io_in(valid_316_io_in),
    .io_out(valid_316_io_out),
    .io_enable(valid_316_io_enable)
  );
  FF_9 valid_317 (
    .clock(valid_317_clock),
    .reset(valid_317_reset),
    .io_in(valid_317_io_in),
    .io_out(valid_317_io_out),
    .io_enable(valid_317_io_enable)
  );
  FF_9 valid_318 (
    .clock(valid_318_clock),
    .reset(valid_318_reset),
    .io_in(valid_318_io_in),
    .io_out(valid_318_io_out),
    .io_enable(valid_318_io_enable)
  );
  FF_9 valid_319 (
    .clock(valid_319_clock),
    .reset(valid_319_reset),
    .io_in(valid_319_io_in),
    .io_out(valid_319_io_out),
    .io_enable(valid_319_io_enable)
  );
  FF_9 valid_320 (
    .clock(valid_320_clock),
    .reset(valid_320_reset),
    .io_in(valid_320_io_in),
    .io_out(valid_320_io_out),
    .io_enable(valid_320_io_enable)
  );
  FF_9 valid_321 (
    .clock(valid_321_clock),
    .reset(valid_321_reset),
    .io_in(valid_321_io_in),
    .io_out(valid_321_io_out),
    .io_enable(valid_321_io_enable)
  );
  FF_9 valid_322 (
    .clock(valid_322_clock),
    .reset(valid_322_reset),
    .io_in(valid_322_io_in),
    .io_out(valid_322_io_out),
    .io_enable(valid_322_io_enable)
  );
  FF_9 valid_323 (
    .clock(valid_323_clock),
    .reset(valid_323_reset),
    .io_in(valid_323_io_in),
    .io_out(valid_323_io_out),
    .io_enable(valid_323_io_enable)
  );
  FF_9 valid_324 (
    .clock(valid_324_clock),
    .reset(valid_324_reset),
    .io_in(valid_324_io_in),
    .io_out(valid_324_io_out),
    .io_enable(valid_324_io_enable)
  );
  FF_9 valid_325 (
    .clock(valid_325_clock),
    .reset(valid_325_reset),
    .io_in(valid_325_io_in),
    .io_out(valid_325_io_out),
    .io_enable(valid_325_io_enable)
  );
  FF_9 valid_326 (
    .clock(valid_326_clock),
    .reset(valid_326_reset),
    .io_in(valid_326_io_in),
    .io_out(valid_326_io_out),
    .io_enable(valid_326_io_enable)
  );
  FF_9 valid_327 (
    .clock(valid_327_clock),
    .reset(valid_327_reset),
    .io_in(valid_327_io_in),
    .io_out(valid_327_io_out),
    .io_enable(valid_327_io_enable)
  );
  FF_9 valid_328 (
    .clock(valid_328_clock),
    .reset(valid_328_reset),
    .io_in(valid_328_io_in),
    .io_out(valid_328_io_out),
    .io_enable(valid_328_io_enable)
  );
  FF_9 valid_329 (
    .clock(valid_329_clock),
    .reset(valid_329_reset),
    .io_in(valid_329_io_in),
    .io_out(valid_329_io_out),
    .io_enable(valid_329_io_enable)
  );
  FF_9 valid_330 (
    .clock(valid_330_clock),
    .reset(valid_330_reset),
    .io_in(valid_330_io_in),
    .io_out(valid_330_io_out),
    .io_enable(valid_330_io_enable)
  );
  FF_9 valid_331 (
    .clock(valid_331_clock),
    .reset(valid_331_reset),
    .io_in(valid_331_io_in),
    .io_out(valid_331_io_out),
    .io_enable(valid_331_io_enable)
  );
  FF_9 valid_332 (
    .clock(valid_332_clock),
    .reset(valid_332_reset),
    .io_in(valid_332_io_in),
    .io_out(valid_332_io_out),
    .io_enable(valid_332_io_enable)
  );
  FF_9 valid_333 (
    .clock(valid_333_clock),
    .reset(valid_333_reset),
    .io_in(valid_333_io_in),
    .io_out(valid_333_io_out),
    .io_enable(valid_333_io_enable)
  );
  FF_9 valid_334 (
    .clock(valid_334_clock),
    .reset(valid_334_reset),
    .io_in(valid_334_io_in),
    .io_out(valid_334_io_out),
    .io_enable(valid_334_io_enable)
  );
  FF_9 valid_335 (
    .clock(valid_335_clock),
    .reset(valid_335_reset),
    .io_in(valid_335_io_in),
    .io_out(valid_335_io_out),
    .io_enable(valid_335_io_enable)
  );
  FF_9 valid_336 (
    .clock(valid_336_clock),
    .reset(valid_336_reset),
    .io_in(valid_336_io_in),
    .io_out(valid_336_io_out),
    .io_enable(valid_336_io_enable)
  );
  FF_9 valid_337 (
    .clock(valid_337_clock),
    .reset(valid_337_reset),
    .io_in(valid_337_io_in),
    .io_out(valid_337_io_out),
    .io_enable(valid_337_io_enable)
  );
  FF_9 valid_338 (
    .clock(valid_338_clock),
    .reset(valid_338_reset),
    .io_in(valid_338_io_in),
    .io_out(valid_338_io_out),
    .io_enable(valid_338_io_enable)
  );
  FF_9 valid_339 (
    .clock(valid_339_clock),
    .reset(valid_339_reset),
    .io_in(valid_339_io_in),
    .io_out(valid_339_io_out),
    .io_enable(valid_339_io_enable)
  );
  FF_9 valid_340 (
    .clock(valid_340_clock),
    .reset(valid_340_reset),
    .io_in(valid_340_io_in),
    .io_out(valid_340_io_out),
    .io_enable(valid_340_io_enable)
  );
  FF_9 valid_341 (
    .clock(valid_341_clock),
    .reset(valid_341_reset),
    .io_in(valid_341_io_in),
    .io_out(valid_341_io_out),
    .io_enable(valid_341_io_enable)
  );
  FF_9 valid_342 (
    .clock(valid_342_clock),
    .reset(valid_342_reset),
    .io_in(valid_342_io_in),
    .io_out(valid_342_io_out),
    .io_enable(valid_342_io_enable)
  );
  FF_9 valid_343 (
    .clock(valid_343_clock),
    .reset(valid_343_reset),
    .io_in(valid_343_io_in),
    .io_out(valid_343_io_out),
    .io_enable(valid_343_io_enable)
  );
  FF_9 valid_344 (
    .clock(valid_344_clock),
    .reset(valid_344_reset),
    .io_in(valid_344_io_in),
    .io_out(valid_344_io_out),
    .io_enable(valid_344_io_enable)
  );
  FF_9 valid_345 (
    .clock(valid_345_clock),
    .reset(valid_345_reset),
    .io_in(valid_345_io_in),
    .io_out(valid_345_io_out),
    .io_enable(valid_345_io_enable)
  );
  FF_9 valid_346 (
    .clock(valid_346_clock),
    .reset(valid_346_reset),
    .io_in(valid_346_io_in),
    .io_out(valid_346_io_out),
    .io_enable(valid_346_io_enable)
  );
  FF_9 valid_347 (
    .clock(valid_347_clock),
    .reset(valid_347_reset),
    .io_in(valid_347_io_in),
    .io_out(valid_347_io_out),
    .io_enable(valid_347_io_enable)
  );
  FF_9 valid_348 (
    .clock(valid_348_clock),
    .reset(valid_348_reset),
    .io_in(valid_348_io_in),
    .io_out(valid_348_io_out),
    .io_enable(valid_348_io_enable)
  );
  FF_9 valid_349 (
    .clock(valid_349_clock),
    .reset(valid_349_reset),
    .io_in(valid_349_io_in),
    .io_out(valid_349_io_out),
    .io_enable(valid_349_io_enable)
  );
  FF_9 valid_350 (
    .clock(valid_350_clock),
    .reset(valid_350_reset),
    .io_in(valid_350_io_in),
    .io_out(valid_350_io_out),
    .io_enable(valid_350_io_enable)
  );
  FF_9 valid_351 (
    .clock(valid_351_clock),
    .reset(valid_351_reset),
    .io_in(valid_351_io_in),
    .io_out(valid_351_io_out),
    .io_enable(valid_351_io_enable)
  );
  FF_9 valid_352 (
    .clock(valid_352_clock),
    .reset(valid_352_reset),
    .io_in(valid_352_io_in),
    .io_out(valid_352_io_out),
    .io_enable(valid_352_io_enable)
  );
  FF_9 valid_353 (
    .clock(valid_353_clock),
    .reset(valid_353_reset),
    .io_in(valid_353_io_in),
    .io_out(valid_353_io_out),
    .io_enable(valid_353_io_enable)
  );
  FF_9 valid_354 (
    .clock(valid_354_clock),
    .reset(valid_354_reset),
    .io_in(valid_354_io_in),
    .io_out(valid_354_io_out),
    .io_enable(valid_354_io_enable)
  );
  FF_9 valid_355 (
    .clock(valid_355_clock),
    .reset(valid_355_reset),
    .io_in(valid_355_io_in),
    .io_out(valid_355_io_out),
    .io_enable(valid_355_io_enable)
  );
  FF_9 valid_356 (
    .clock(valid_356_clock),
    .reset(valid_356_reset),
    .io_in(valid_356_io_in),
    .io_out(valid_356_io_out),
    .io_enable(valid_356_io_enable)
  );
  FF_9 valid_357 (
    .clock(valid_357_clock),
    .reset(valid_357_reset),
    .io_in(valid_357_io_in),
    .io_out(valid_357_io_out),
    .io_enable(valid_357_io_enable)
  );
  FF_9 valid_358 (
    .clock(valid_358_clock),
    .reset(valid_358_reset),
    .io_in(valid_358_io_in),
    .io_out(valid_358_io_out),
    .io_enable(valid_358_io_enable)
  );
  FF_9 valid_359 (
    .clock(valid_359_clock),
    .reset(valid_359_reset),
    .io_in(valid_359_io_in),
    .io_out(valid_359_io_out),
    .io_enable(valid_359_io_enable)
  );
  FF_9 valid_360 (
    .clock(valid_360_clock),
    .reset(valid_360_reset),
    .io_in(valid_360_io_in),
    .io_out(valid_360_io_out),
    .io_enable(valid_360_io_enable)
  );
  FF_9 valid_361 (
    .clock(valid_361_clock),
    .reset(valid_361_reset),
    .io_in(valid_361_io_in),
    .io_out(valid_361_io_out),
    .io_enable(valid_361_io_enable)
  );
  FF_9 valid_362 (
    .clock(valid_362_clock),
    .reset(valid_362_reset),
    .io_in(valid_362_io_in),
    .io_out(valid_362_io_out),
    .io_enable(valid_362_io_enable)
  );
  FF_9 valid_363 (
    .clock(valid_363_clock),
    .reset(valid_363_reset),
    .io_in(valid_363_io_in),
    .io_out(valid_363_io_out),
    .io_enable(valid_363_io_enable)
  );
  FF_9 valid_364 (
    .clock(valid_364_clock),
    .reset(valid_364_reset),
    .io_in(valid_364_io_in),
    .io_out(valid_364_io_out),
    .io_enable(valid_364_io_enable)
  );
  FF_9 valid_365 (
    .clock(valid_365_clock),
    .reset(valid_365_reset),
    .io_in(valid_365_io_in),
    .io_out(valid_365_io_out),
    .io_enable(valid_365_io_enable)
  );
  FF_9 valid_366 (
    .clock(valid_366_clock),
    .reset(valid_366_reset),
    .io_in(valid_366_io_in),
    .io_out(valid_366_io_out),
    .io_enable(valid_366_io_enable)
  );
  FF_9 valid_367 (
    .clock(valid_367_clock),
    .reset(valid_367_reset),
    .io_in(valid_367_io_in),
    .io_out(valid_367_io_out),
    .io_enable(valid_367_io_enable)
  );
  FF_9 valid_368 (
    .clock(valid_368_clock),
    .reset(valid_368_reset),
    .io_in(valid_368_io_in),
    .io_out(valid_368_io_out),
    .io_enable(valid_368_io_enable)
  );
  FF_9 valid_369 (
    .clock(valid_369_clock),
    .reset(valid_369_reset),
    .io_in(valid_369_io_in),
    .io_out(valid_369_io_out),
    .io_enable(valid_369_io_enable)
  );
  FF_9 valid_370 (
    .clock(valid_370_clock),
    .reset(valid_370_reset),
    .io_in(valid_370_io_in),
    .io_out(valid_370_io_out),
    .io_enable(valid_370_io_enable)
  );
  FF_9 valid_371 (
    .clock(valid_371_clock),
    .reset(valid_371_reset),
    .io_in(valid_371_io_in),
    .io_out(valid_371_io_out),
    .io_enable(valid_371_io_enable)
  );
  FF_9 valid_372 (
    .clock(valid_372_clock),
    .reset(valid_372_reset),
    .io_in(valid_372_io_in),
    .io_out(valid_372_io_out),
    .io_enable(valid_372_io_enable)
  );
  FF_9 valid_373 (
    .clock(valid_373_clock),
    .reset(valid_373_reset),
    .io_in(valid_373_io_in),
    .io_out(valid_373_io_out),
    .io_enable(valid_373_io_enable)
  );
  FF_9 valid_374 (
    .clock(valid_374_clock),
    .reset(valid_374_reset),
    .io_in(valid_374_io_in),
    .io_out(valid_374_io_out),
    .io_enable(valid_374_io_enable)
  );
  FF_9 valid_375 (
    .clock(valid_375_clock),
    .reset(valid_375_reset),
    .io_in(valid_375_io_in),
    .io_out(valid_375_io_out),
    .io_enable(valid_375_io_enable)
  );
  FF_9 valid_376 (
    .clock(valid_376_clock),
    .reset(valid_376_reset),
    .io_in(valid_376_io_in),
    .io_out(valid_376_io_out),
    .io_enable(valid_376_io_enable)
  );
  FF_9 valid_377 (
    .clock(valid_377_clock),
    .reset(valid_377_reset),
    .io_in(valid_377_io_in),
    .io_out(valid_377_io_out),
    .io_enable(valid_377_io_enable)
  );
  FF_9 valid_378 (
    .clock(valid_378_clock),
    .reset(valid_378_reset),
    .io_in(valid_378_io_in),
    .io_out(valid_378_io_out),
    .io_enable(valid_378_io_enable)
  );
  FF_9 valid_379 (
    .clock(valid_379_clock),
    .reset(valid_379_reset),
    .io_in(valid_379_io_in),
    .io_out(valid_379_io_out),
    .io_enable(valid_379_io_enable)
  );
  FF_9 valid_380 (
    .clock(valid_380_clock),
    .reset(valid_380_reset),
    .io_in(valid_380_io_in),
    .io_out(valid_380_io_out),
    .io_enable(valid_380_io_enable)
  );
  FF_9 valid_381 (
    .clock(valid_381_clock),
    .reset(valid_381_reset),
    .io_in(valid_381_io_in),
    .io_out(valid_381_io_out),
    .io_enable(valid_381_io_enable)
  );
  FF_9 valid_382 (
    .clock(valid_382_clock),
    .reset(valid_382_reset),
    .io_in(valid_382_io_in),
    .io_out(valid_382_io_out),
    .io_enable(valid_382_io_enable)
  );
  FF_9 valid_383 (
    .clock(valid_383_clock),
    .reset(valid_383_reset),
    .io_in(valid_383_io_in),
    .io_out(valid_383_io_out),
    .io_enable(valid_383_io_enable)
  );
  FF_9 valid_384 (
    .clock(valid_384_clock),
    .reset(valid_384_reset),
    .io_in(valid_384_io_in),
    .io_out(valid_384_io_out),
    .io_enable(valid_384_io_enable)
  );
  FF_9 valid_385 (
    .clock(valid_385_clock),
    .reset(valid_385_reset),
    .io_in(valid_385_io_in),
    .io_out(valid_385_io_out),
    .io_enable(valid_385_io_enable)
  );
  FF_9 valid_386 (
    .clock(valid_386_clock),
    .reset(valid_386_reset),
    .io_in(valid_386_io_in),
    .io_out(valid_386_io_out),
    .io_enable(valid_386_io_enable)
  );
  FF_9 valid_387 (
    .clock(valid_387_clock),
    .reset(valid_387_reset),
    .io_in(valid_387_io_in),
    .io_out(valid_387_io_out),
    .io_enable(valid_387_io_enable)
  );
  FF_9 valid_388 (
    .clock(valid_388_clock),
    .reset(valid_388_reset),
    .io_in(valid_388_io_in),
    .io_out(valid_388_io_out),
    .io_enable(valid_388_io_enable)
  );
  FF_9 valid_389 (
    .clock(valid_389_clock),
    .reset(valid_389_reset),
    .io_in(valid_389_io_in),
    .io_out(valid_389_io_out),
    .io_enable(valid_389_io_enable)
  );
  FF_9 valid_390 (
    .clock(valid_390_clock),
    .reset(valid_390_reset),
    .io_in(valid_390_io_in),
    .io_out(valid_390_io_out),
    .io_enable(valid_390_io_enable)
  );
  FF_9 valid_391 (
    .clock(valid_391_clock),
    .reset(valid_391_reset),
    .io_in(valid_391_io_in),
    .io_out(valid_391_io_out),
    .io_enable(valid_391_io_enable)
  );
  FF_9 valid_392 (
    .clock(valid_392_clock),
    .reset(valid_392_reset),
    .io_in(valid_392_io_in),
    .io_out(valid_392_io_out),
    .io_enable(valid_392_io_enable)
  );
  FF_9 valid_393 (
    .clock(valid_393_clock),
    .reset(valid_393_reset),
    .io_in(valid_393_io_in),
    .io_out(valid_393_io_out),
    .io_enable(valid_393_io_enable)
  );
  FF_9 valid_394 (
    .clock(valid_394_clock),
    .reset(valid_394_reset),
    .io_in(valid_394_io_in),
    .io_out(valid_394_io_out),
    .io_enable(valid_394_io_enable)
  );
  FF_9 valid_395 (
    .clock(valid_395_clock),
    .reset(valid_395_reset),
    .io_in(valid_395_io_in),
    .io_out(valid_395_io_out),
    .io_enable(valid_395_io_enable)
  );
  FF_9 valid_396 (
    .clock(valid_396_clock),
    .reset(valid_396_reset),
    .io_in(valid_396_io_in),
    .io_out(valid_396_io_out),
    .io_enable(valid_396_io_enable)
  );
  FF_9 valid_397 (
    .clock(valid_397_clock),
    .reset(valid_397_reset),
    .io_in(valid_397_io_in),
    .io_out(valid_397_io_out),
    .io_enable(valid_397_io_enable)
  );
  FF_9 valid_398 (
    .clock(valid_398_clock),
    .reset(valid_398_reset),
    .io_in(valid_398_io_in),
    .io_out(valid_398_io_out),
    .io_enable(valid_398_io_enable)
  );
  FF_9 valid_399 (
    .clock(valid_399_clock),
    .reset(valid_399_reset),
    .io_in(valid_399_io_in),
    .io_out(valid_399_io_out),
    .io_enable(valid_399_io_enable)
  );
  FF_9 valid_400 (
    .clock(valid_400_clock),
    .reset(valid_400_reset),
    .io_in(valid_400_io_in),
    .io_out(valid_400_io_out),
    .io_enable(valid_400_io_enable)
  );
  FF_9 valid_401 (
    .clock(valid_401_clock),
    .reset(valid_401_reset),
    .io_in(valid_401_io_in),
    .io_out(valid_401_io_out),
    .io_enable(valid_401_io_enable)
  );
  FF_9 valid_402 (
    .clock(valid_402_clock),
    .reset(valid_402_reset),
    .io_in(valid_402_io_in),
    .io_out(valid_402_io_out),
    .io_enable(valid_402_io_enable)
  );
  FF_9 valid_403 (
    .clock(valid_403_clock),
    .reset(valid_403_reset),
    .io_in(valid_403_io_in),
    .io_out(valid_403_io_out),
    .io_enable(valid_403_io_enable)
  );
  FF_9 valid_404 (
    .clock(valid_404_clock),
    .reset(valid_404_reset),
    .io_in(valid_404_io_in),
    .io_out(valid_404_io_out),
    .io_enable(valid_404_io_enable)
  );
  FF_9 valid_405 (
    .clock(valid_405_clock),
    .reset(valid_405_reset),
    .io_in(valid_405_io_in),
    .io_out(valid_405_io_out),
    .io_enable(valid_405_io_enable)
  );
  FF_9 valid_406 (
    .clock(valid_406_clock),
    .reset(valid_406_reset),
    .io_in(valid_406_io_in),
    .io_out(valid_406_io_out),
    .io_enable(valid_406_io_enable)
  );
  FF_9 valid_407 (
    .clock(valid_407_clock),
    .reset(valid_407_reset),
    .io_in(valid_407_io_in),
    .io_out(valid_407_io_out),
    .io_enable(valid_407_io_enable)
  );
  FF_9 valid_408 (
    .clock(valid_408_clock),
    .reset(valid_408_reset),
    .io_in(valid_408_io_in),
    .io_out(valid_408_io_out),
    .io_enable(valid_408_io_enable)
  );
  FF_9 valid_409 (
    .clock(valid_409_clock),
    .reset(valid_409_reset),
    .io_in(valid_409_io_in),
    .io_out(valid_409_io_out),
    .io_enable(valid_409_io_enable)
  );
  FF_9 valid_410 (
    .clock(valid_410_clock),
    .reset(valid_410_reset),
    .io_in(valid_410_io_in),
    .io_out(valid_410_io_out),
    .io_enable(valid_410_io_enable)
  );
  FF_9 valid_411 (
    .clock(valid_411_clock),
    .reset(valid_411_reset),
    .io_in(valid_411_io_in),
    .io_out(valid_411_io_out),
    .io_enable(valid_411_io_enable)
  );
  FF_9 valid_412 (
    .clock(valid_412_clock),
    .reset(valid_412_reset),
    .io_in(valid_412_io_in),
    .io_out(valid_412_io_out),
    .io_enable(valid_412_io_enable)
  );
  FF_9 valid_413 (
    .clock(valid_413_clock),
    .reset(valid_413_reset),
    .io_in(valid_413_io_in),
    .io_out(valid_413_io_out),
    .io_enable(valid_413_io_enable)
  );
  FF_9 valid_414 (
    .clock(valid_414_clock),
    .reset(valid_414_reset),
    .io_in(valid_414_io_in),
    .io_out(valid_414_io_out),
    .io_enable(valid_414_io_enable)
  );
  FF_9 valid_415 (
    .clock(valid_415_clock),
    .reset(valid_415_reset),
    .io_in(valid_415_io_in),
    .io_out(valid_415_io_out),
    .io_enable(valid_415_io_enable)
  );
  FF_9 valid_416 (
    .clock(valid_416_clock),
    .reset(valid_416_reset),
    .io_in(valid_416_io_in),
    .io_out(valid_416_io_out),
    .io_enable(valid_416_io_enable)
  );
  FF_9 valid_417 (
    .clock(valid_417_clock),
    .reset(valid_417_reset),
    .io_in(valid_417_io_in),
    .io_out(valid_417_io_out),
    .io_enable(valid_417_io_enable)
  );
  FF_9 valid_418 (
    .clock(valid_418_clock),
    .reset(valid_418_reset),
    .io_in(valid_418_io_in),
    .io_out(valid_418_io_out),
    .io_enable(valid_418_io_enable)
  );
  FF_9 valid_419 (
    .clock(valid_419_clock),
    .reset(valid_419_reset),
    .io_in(valid_419_io_in),
    .io_out(valid_419_io_out),
    .io_enable(valid_419_io_enable)
  );
  FF_9 valid_420 (
    .clock(valid_420_clock),
    .reset(valid_420_reset),
    .io_in(valid_420_io_in),
    .io_out(valid_420_io_out),
    .io_enable(valid_420_io_enable)
  );
  FF_9 valid_421 (
    .clock(valid_421_clock),
    .reset(valid_421_reset),
    .io_in(valid_421_io_in),
    .io_out(valid_421_io_out),
    .io_enable(valid_421_io_enable)
  );
  FF_9 valid_422 (
    .clock(valid_422_clock),
    .reset(valid_422_reset),
    .io_in(valid_422_io_in),
    .io_out(valid_422_io_out),
    .io_enable(valid_422_io_enable)
  );
  FF_9 valid_423 (
    .clock(valid_423_clock),
    .reset(valid_423_reset),
    .io_in(valid_423_io_in),
    .io_out(valid_423_io_out),
    .io_enable(valid_423_io_enable)
  );
  FF_9 valid_424 (
    .clock(valid_424_clock),
    .reset(valid_424_reset),
    .io_in(valid_424_io_in),
    .io_out(valid_424_io_out),
    .io_enable(valid_424_io_enable)
  );
  FF_9 valid_425 (
    .clock(valid_425_clock),
    .reset(valid_425_reset),
    .io_in(valid_425_io_in),
    .io_out(valid_425_io_out),
    .io_enable(valid_425_io_enable)
  );
  FF_9 valid_426 (
    .clock(valid_426_clock),
    .reset(valid_426_reset),
    .io_in(valid_426_io_in),
    .io_out(valid_426_io_out),
    .io_enable(valid_426_io_enable)
  );
  FF_9 valid_427 (
    .clock(valid_427_clock),
    .reset(valid_427_reset),
    .io_in(valid_427_io_in),
    .io_out(valid_427_io_out),
    .io_enable(valid_427_io_enable)
  );
  FF_9 valid_428 (
    .clock(valid_428_clock),
    .reset(valid_428_reset),
    .io_in(valid_428_io_in),
    .io_out(valid_428_io_out),
    .io_enable(valid_428_io_enable)
  );
  FF_9 valid_429 (
    .clock(valid_429_clock),
    .reset(valid_429_reset),
    .io_in(valid_429_io_in),
    .io_out(valid_429_io_out),
    .io_enable(valid_429_io_enable)
  );
  FF_9 valid_430 (
    .clock(valid_430_clock),
    .reset(valid_430_reset),
    .io_in(valid_430_io_in),
    .io_out(valid_430_io_out),
    .io_enable(valid_430_io_enable)
  );
  FF_9 valid_431 (
    .clock(valid_431_clock),
    .reset(valid_431_reset),
    .io_in(valid_431_io_in),
    .io_out(valid_431_io_out),
    .io_enable(valid_431_io_enable)
  );
  FF_9 valid_432 (
    .clock(valid_432_clock),
    .reset(valid_432_reset),
    .io_in(valid_432_io_in),
    .io_out(valid_432_io_out),
    .io_enable(valid_432_io_enable)
  );
  FF_9 valid_433 (
    .clock(valid_433_clock),
    .reset(valid_433_reset),
    .io_in(valid_433_io_in),
    .io_out(valid_433_io_out),
    .io_enable(valid_433_io_enable)
  );
  FF_9 valid_434 (
    .clock(valid_434_clock),
    .reset(valid_434_reset),
    .io_in(valid_434_io_in),
    .io_out(valid_434_io_out),
    .io_enable(valid_434_io_enable)
  );
  FF_9 valid_435 (
    .clock(valid_435_clock),
    .reset(valid_435_reset),
    .io_in(valid_435_io_in),
    .io_out(valid_435_io_out),
    .io_enable(valid_435_io_enable)
  );
  FF_9 valid_436 (
    .clock(valid_436_clock),
    .reset(valid_436_reset),
    .io_in(valid_436_io_in),
    .io_out(valid_436_io_out),
    .io_enable(valid_436_io_enable)
  );
  FF_9 valid_437 (
    .clock(valid_437_clock),
    .reset(valid_437_reset),
    .io_in(valid_437_io_in),
    .io_out(valid_437_io_out),
    .io_enable(valid_437_io_enable)
  );
  FF_9 valid_438 (
    .clock(valid_438_clock),
    .reset(valid_438_reset),
    .io_in(valid_438_io_in),
    .io_out(valid_438_io_out),
    .io_enable(valid_438_io_enable)
  );
  FF_9 valid_439 (
    .clock(valid_439_clock),
    .reset(valid_439_reset),
    .io_in(valid_439_io_in),
    .io_out(valid_439_io_out),
    .io_enable(valid_439_io_enable)
  );
  FF_9 valid_440 (
    .clock(valid_440_clock),
    .reset(valid_440_reset),
    .io_in(valid_440_io_in),
    .io_out(valid_440_io_out),
    .io_enable(valid_440_io_enable)
  );
  FF_9 valid_441 (
    .clock(valid_441_clock),
    .reset(valid_441_reset),
    .io_in(valid_441_io_in),
    .io_out(valid_441_io_out),
    .io_enable(valid_441_io_enable)
  );
  FF_9 valid_442 (
    .clock(valid_442_clock),
    .reset(valid_442_reset),
    .io_in(valid_442_io_in),
    .io_out(valid_442_io_out),
    .io_enable(valid_442_io_enable)
  );
  FF_9 valid_443 (
    .clock(valid_443_clock),
    .reset(valid_443_reset),
    .io_in(valid_443_io_in),
    .io_out(valid_443_io_out),
    .io_enable(valid_443_io_enable)
  );
  FF_9 valid_444 (
    .clock(valid_444_clock),
    .reset(valid_444_reset),
    .io_in(valid_444_io_in),
    .io_out(valid_444_io_out),
    .io_enable(valid_444_io_enable)
  );
  FF_9 valid_445 (
    .clock(valid_445_clock),
    .reset(valid_445_reset),
    .io_in(valid_445_io_in),
    .io_out(valid_445_io_out),
    .io_enable(valid_445_io_enable)
  );
  FF_9 valid_446 (
    .clock(valid_446_clock),
    .reset(valid_446_reset),
    .io_in(valid_446_io_in),
    .io_out(valid_446_io_out),
    .io_enable(valid_446_io_enable)
  );
  FF_9 valid_447 (
    .clock(valid_447_clock),
    .reset(valid_447_reset),
    .io_in(valid_447_io_in),
    .io_out(valid_447_io_out),
    .io_enable(valid_447_io_enable)
  );
  FF_9 valid_448 (
    .clock(valid_448_clock),
    .reset(valid_448_reset),
    .io_in(valid_448_io_in),
    .io_out(valid_448_io_out),
    .io_enable(valid_448_io_enable)
  );
  FF_9 valid_449 (
    .clock(valid_449_clock),
    .reset(valid_449_reset),
    .io_in(valid_449_io_in),
    .io_out(valid_449_io_out),
    .io_enable(valid_449_io_enable)
  );
  FF_9 valid_450 (
    .clock(valid_450_clock),
    .reset(valid_450_reset),
    .io_in(valid_450_io_in),
    .io_out(valid_450_io_out),
    .io_enable(valid_450_io_enable)
  );
  FF_9 valid_451 (
    .clock(valid_451_clock),
    .reset(valid_451_reset),
    .io_in(valid_451_io_in),
    .io_out(valid_451_io_out),
    .io_enable(valid_451_io_enable)
  );
  FF_9 valid_452 (
    .clock(valid_452_clock),
    .reset(valid_452_reset),
    .io_in(valid_452_io_in),
    .io_out(valid_452_io_out),
    .io_enable(valid_452_io_enable)
  );
  FF_9 valid_453 (
    .clock(valid_453_clock),
    .reset(valid_453_reset),
    .io_in(valid_453_io_in),
    .io_out(valid_453_io_out),
    .io_enable(valid_453_io_enable)
  );
  FF_9 valid_454 (
    .clock(valid_454_clock),
    .reset(valid_454_reset),
    .io_in(valid_454_io_in),
    .io_out(valid_454_io_out),
    .io_enable(valid_454_io_enable)
  );
  FF_9 valid_455 (
    .clock(valid_455_clock),
    .reset(valid_455_reset),
    .io_in(valid_455_io_in),
    .io_out(valid_455_io_out),
    .io_enable(valid_455_io_enable)
  );
  FF_9 valid_456 (
    .clock(valid_456_clock),
    .reset(valid_456_reset),
    .io_in(valid_456_io_in),
    .io_out(valid_456_io_out),
    .io_enable(valid_456_io_enable)
  );
  FF_9 valid_457 (
    .clock(valid_457_clock),
    .reset(valid_457_reset),
    .io_in(valid_457_io_in),
    .io_out(valid_457_io_out),
    .io_enable(valid_457_io_enable)
  );
  FF_9 valid_458 (
    .clock(valid_458_clock),
    .reset(valid_458_reset),
    .io_in(valid_458_io_in),
    .io_out(valid_458_io_out),
    .io_enable(valid_458_io_enable)
  );
  FF_9 valid_459 (
    .clock(valid_459_clock),
    .reset(valid_459_reset),
    .io_in(valid_459_io_in),
    .io_out(valid_459_io_out),
    .io_enable(valid_459_io_enable)
  );
  FF_9 valid_460 (
    .clock(valid_460_clock),
    .reset(valid_460_reset),
    .io_in(valid_460_io_in),
    .io_out(valid_460_io_out),
    .io_enable(valid_460_io_enable)
  );
  FF_9 valid_461 (
    .clock(valid_461_clock),
    .reset(valid_461_reset),
    .io_in(valid_461_io_in),
    .io_out(valid_461_io_out),
    .io_enable(valid_461_io_enable)
  );
  FF_9 valid_462 (
    .clock(valid_462_clock),
    .reset(valid_462_reset),
    .io_in(valid_462_io_in),
    .io_out(valid_462_io_out),
    .io_enable(valid_462_io_enable)
  );
  FF_9 valid_463 (
    .clock(valid_463_clock),
    .reset(valid_463_reset),
    .io_in(valid_463_io_in),
    .io_out(valid_463_io_out),
    .io_enable(valid_463_io_enable)
  );
  FF_9 valid_464 (
    .clock(valid_464_clock),
    .reset(valid_464_reset),
    .io_in(valid_464_io_in),
    .io_out(valid_464_io_out),
    .io_enable(valid_464_io_enable)
  );
  FF_9 valid_465 (
    .clock(valid_465_clock),
    .reset(valid_465_reset),
    .io_in(valid_465_io_in),
    .io_out(valid_465_io_out),
    .io_enable(valid_465_io_enable)
  );
  FF_9 valid_466 (
    .clock(valid_466_clock),
    .reset(valid_466_reset),
    .io_in(valid_466_io_in),
    .io_out(valid_466_io_out),
    .io_enable(valid_466_io_enable)
  );
  FF_9 valid_467 (
    .clock(valid_467_clock),
    .reset(valid_467_reset),
    .io_in(valid_467_io_in),
    .io_out(valid_467_io_out),
    .io_enable(valid_467_io_enable)
  );
  FF_9 valid_468 (
    .clock(valid_468_clock),
    .reset(valid_468_reset),
    .io_in(valid_468_io_in),
    .io_out(valid_468_io_out),
    .io_enable(valid_468_io_enable)
  );
  FF_9 valid_469 (
    .clock(valid_469_clock),
    .reset(valid_469_reset),
    .io_in(valid_469_io_in),
    .io_out(valid_469_io_out),
    .io_enable(valid_469_io_enable)
  );
  FF_9 valid_470 (
    .clock(valid_470_clock),
    .reset(valid_470_reset),
    .io_in(valid_470_io_in),
    .io_out(valid_470_io_out),
    .io_enable(valid_470_io_enable)
  );
  FF_9 valid_471 (
    .clock(valid_471_clock),
    .reset(valid_471_reset),
    .io_in(valid_471_io_in),
    .io_out(valid_471_io_out),
    .io_enable(valid_471_io_enable)
  );
  FF_9 valid_472 (
    .clock(valid_472_clock),
    .reset(valid_472_reset),
    .io_in(valid_472_io_in),
    .io_out(valid_472_io_out),
    .io_enable(valid_472_io_enable)
  );
  FF_9 valid_473 (
    .clock(valid_473_clock),
    .reset(valid_473_reset),
    .io_in(valid_473_io_in),
    .io_out(valid_473_io_out),
    .io_enable(valid_473_io_enable)
  );
  FF_9 valid_474 (
    .clock(valid_474_clock),
    .reset(valid_474_reset),
    .io_in(valid_474_io_in),
    .io_out(valid_474_io_out),
    .io_enable(valid_474_io_enable)
  );
  FF_9 valid_475 (
    .clock(valid_475_clock),
    .reset(valid_475_reset),
    .io_in(valid_475_io_in),
    .io_out(valid_475_io_out),
    .io_enable(valid_475_io_enable)
  );
  FF_9 valid_476 (
    .clock(valid_476_clock),
    .reset(valid_476_reset),
    .io_in(valid_476_io_in),
    .io_out(valid_476_io_out),
    .io_enable(valid_476_io_enable)
  );
  FF_9 valid_477 (
    .clock(valid_477_clock),
    .reset(valid_477_reset),
    .io_in(valid_477_io_in),
    .io_out(valid_477_io_out),
    .io_enable(valid_477_io_enable)
  );
  FF_9 valid_478 (
    .clock(valid_478_clock),
    .reset(valid_478_reset),
    .io_in(valid_478_io_in),
    .io_out(valid_478_io_out),
    .io_enable(valid_478_io_enable)
  );
  FF_9 valid_479 (
    .clock(valid_479_clock),
    .reset(valid_479_reset),
    .io_in(valid_479_io_in),
    .io_out(valid_479_io_out),
    .io_enable(valid_479_io_enable)
  );
  FF_9 valid_480 (
    .clock(valid_480_clock),
    .reset(valid_480_reset),
    .io_in(valid_480_io_in),
    .io_out(valid_480_io_out),
    .io_enable(valid_480_io_enable)
  );
  FF_9 valid_481 (
    .clock(valid_481_clock),
    .reset(valid_481_reset),
    .io_in(valid_481_io_in),
    .io_out(valid_481_io_out),
    .io_enable(valid_481_io_enable)
  );
  FF_9 valid_482 (
    .clock(valid_482_clock),
    .reset(valid_482_reset),
    .io_in(valid_482_io_in),
    .io_out(valid_482_io_out),
    .io_enable(valid_482_io_enable)
  );
  FF_9 valid_483 (
    .clock(valid_483_clock),
    .reset(valid_483_reset),
    .io_in(valid_483_io_in),
    .io_out(valid_483_io_out),
    .io_enable(valid_483_io_enable)
  );
  FF_9 valid_484 (
    .clock(valid_484_clock),
    .reset(valid_484_reset),
    .io_in(valid_484_io_in),
    .io_out(valid_484_io_out),
    .io_enable(valid_484_io_enable)
  );
  FF_9 valid_485 (
    .clock(valid_485_clock),
    .reset(valid_485_reset),
    .io_in(valid_485_io_in),
    .io_out(valid_485_io_out),
    .io_enable(valid_485_io_enable)
  );
  FF_9 valid_486 (
    .clock(valid_486_clock),
    .reset(valid_486_reset),
    .io_in(valid_486_io_in),
    .io_out(valid_486_io_out),
    .io_enable(valid_486_io_enable)
  );
  FF_9 valid_487 (
    .clock(valid_487_clock),
    .reset(valid_487_reset),
    .io_in(valid_487_io_in),
    .io_out(valid_487_io_out),
    .io_enable(valid_487_io_enable)
  );
  FF_9 valid_488 (
    .clock(valid_488_clock),
    .reset(valid_488_reset),
    .io_in(valid_488_io_in),
    .io_out(valid_488_io_out),
    .io_enable(valid_488_io_enable)
  );
  FF_9 valid_489 (
    .clock(valid_489_clock),
    .reset(valid_489_reset),
    .io_in(valid_489_io_in),
    .io_out(valid_489_io_out),
    .io_enable(valid_489_io_enable)
  );
  FF_9 valid_490 (
    .clock(valid_490_clock),
    .reset(valid_490_reset),
    .io_in(valid_490_io_in),
    .io_out(valid_490_io_out),
    .io_enable(valid_490_io_enable)
  );
  FF_9 valid_491 (
    .clock(valid_491_clock),
    .reset(valid_491_reset),
    .io_in(valid_491_io_in),
    .io_out(valid_491_io_out),
    .io_enable(valid_491_io_enable)
  );
  FF_9 valid_492 (
    .clock(valid_492_clock),
    .reset(valid_492_reset),
    .io_in(valid_492_io_in),
    .io_out(valid_492_io_out),
    .io_enable(valid_492_io_enable)
  );
  FF_9 valid_493 (
    .clock(valid_493_clock),
    .reset(valid_493_reset),
    .io_in(valid_493_io_in),
    .io_out(valid_493_io_out),
    .io_enable(valid_493_io_enable)
  );
  FF_9 valid_494 (
    .clock(valid_494_clock),
    .reset(valid_494_reset),
    .io_in(valid_494_io_in),
    .io_out(valid_494_io_out),
    .io_enable(valid_494_io_enable)
  );
  FF_9 valid_495 (
    .clock(valid_495_clock),
    .reset(valid_495_reset),
    .io_in(valid_495_io_in),
    .io_out(valid_495_io_out),
    .io_enable(valid_495_io_enable)
  );
  FF_9 valid_496 (
    .clock(valid_496_clock),
    .reset(valid_496_reset),
    .io_in(valid_496_io_in),
    .io_out(valid_496_io_out),
    .io_enable(valid_496_io_enable)
  );
  FF_9 valid_497 (
    .clock(valid_497_clock),
    .reset(valid_497_reset),
    .io_in(valid_497_io_in),
    .io_out(valid_497_io_out),
    .io_enable(valid_497_io_enable)
  );
  FF_9 valid_498 (
    .clock(valid_498_clock),
    .reset(valid_498_reset),
    .io_in(valid_498_io_in),
    .io_out(valid_498_io_out),
    .io_enable(valid_498_io_enable)
  );
  FF_9 valid_499 (
    .clock(valid_499_clock),
    .reset(valid_499_reset),
    .io_in(valid_499_io_in),
    .io_out(valid_499_io_out),
    .io_enable(valid_499_io_enable)
  );
  FF_9 valid_500 (
    .clock(valid_500_clock),
    .reset(valid_500_reset),
    .io_in(valid_500_io_in),
    .io_out(valid_500_io_out),
    .io_enable(valid_500_io_enable)
  );
  FF_9 valid_501 (
    .clock(valid_501_clock),
    .reset(valid_501_reset),
    .io_in(valid_501_io_in),
    .io_out(valid_501_io_out),
    .io_enable(valid_501_io_enable)
  );
  FF_9 valid_502 (
    .clock(valid_502_clock),
    .reset(valid_502_reset),
    .io_in(valid_502_io_in),
    .io_out(valid_502_io_out),
    .io_enable(valid_502_io_enable)
  );
  FF_9 valid_503 (
    .clock(valid_503_clock),
    .reset(valid_503_reset),
    .io_in(valid_503_io_in),
    .io_out(valid_503_io_out),
    .io_enable(valid_503_io_enable)
  );
  FF_9 valid_504 (
    .clock(valid_504_clock),
    .reset(valid_504_reset),
    .io_in(valid_504_io_in),
    .io_out(valid_504_io_out),
    .io_enable(valid_504_io_enable)
  );
  FF_9 valid_505 (
    .clock(valid_505_clock),
    .reset(valid_505_reset),
    .io_in(valid_505_io_in),
    .io_out(valid_505_io_out),
    .io_enable(valid_505_io_enable)
  );
  FF_9 valid_506 (
    .clock(valid_506_clock),
    .reset(valid_506_reset),
    .io_in(valid_506_io_in),
    .io_out(valid_506_io_out),
    .io_enable(valid_506_io_enable)
  );
  FF_9 valid_507 (
    .clock(valid_507_clock),
    .reset(valid_507_reset),
    .io_in(valid_507_io_in),
    .io_out(valid_507_io_out),
    .io_enable(valid_507_io_enable)
  );
  FF_9 valid_508 (
    .clock(valid_508_clock),
    .reset(valid_508_reset),
    .io_in(valid_508_io_in),
    .io_out(valid_508_io_out),
    .io_enable(valid_508_io_enable)
  );
  FF_9 valid_509 (
    .clock(valid_509_clock),
    .reset(valid_509_reset),
    .io_in(valid_509_io_in),
    .io_out(valid_509_io_out),
    .io_enable(valid_509_io_enable)
  );
  FF_9 valid_510 (
    .clock(valid_510_clock),
    .reset(valid_510_reset),
    .io_in(valid_510_io_in),
    .io_out(valid_510_io_out),
    .io_enable(valid_510_io_enable)
  );
  FF_9 valid_511 (
    .clock(valid_511_clock),
    .reset(valid_511_reset),
    .io_in(valid_511_io_in),
    .io_out(valid_511_io_out),
    .io_enable(valid_511_io_enable)
  );
  FF_558 tags_0 (
    .clock(tags_0_clock),
    .reset(tags_0_reset)
  );
  FF_558 tags_1 (
    .clock(tags_1_clock),
    .reset(tags_1_reset)
  );
  FF_558 tags_2 (
    .clock(tags_2_clock),
    .reset(tags_2_reset)
  );
  FF_558 tags_3 (
    .clock(tags_3_clock),
    .reset(tags_3_reset)
  );
  FF_558 tags_4 (
    .clock(tags_4_clock),
    .reset(tags_4_reset)
  );
  FF_558 tags_5 (
    .clock(tags_5_clock),
    .reset(tags_5_reset)
  );
  FF_558 tags_6 (
    .clock(tags_6_clock),
    .reset(tags_6_reset)
  );
  FF_558 tags_7 (
    .clock(tags_7_clock),
    .reset(tags_7_reset)
  );
  FF_558 tags_8 (
    .clock(tags_8_clock),
    .reset(tags_8_reset)
  );
  FF_558 tags_9 (
    .clock(tags_9_clock),
    .reset(tags_9_reset)
  );
  FF_558 tags_10 (
    .clock(tags_10_clock),
    .reset(tags_10_reset)
  );
  FF_558 tags_11 (
    .clock(tags_11_clock),
    .reset(tags_11_reset)
  );
  FF_558 tags_12 (
    .clock(tags_12_clock),
    .reset(tags_12_reset)
  );
  FF_558 tags_13 (
    .clock(tags_13_clock),
    .reset(tags_13_reset)
  );
  FF_558 tags_14 (
    .clock(tags_14_clock),
    .reset(tags_14_reset)
  );
  FF_558 tags_15 (
    .clock(tags_15_clock),
    .reset(tags_15_reset)
  );
  FF_558 tags_16 (
    .clock(tags_16_clock),
    .reset(tags_16_reset)
  );
  FF_558 tags_17 (
    .clock(tags_17_clock),
    .reset(tags_17_reset)
  );
  FF_558 tags_18 (
    .clock(tags_18_clock),
    .reset(tags_18_reset)
  );
  FF_558 tags_19 (
    .clock(tags_19_clock),
    .reset(tags_19_reset)
  );
  FF_558 tags_20 (
    .clock(tags_20_clock),
    .reset(tags_20_reset)
  );
  FF_558 tags_21 (
    .clock(tags_21_clock),
    .reset(tags_21_reset)
  );
  FF_558 tags_22 (
    .clock(tags_22_clock),
    .reset(tags_22_reset)
  );
  FF_558 tags_23 (
    .clock(tags_23_clock),
    .reset(tags_23_reset)
  );
  FF_558 tags_24 (
    .clock(tags_24_clock),
    .reset(tags_24_reset)
  );
  FF_558 tags_25 (
    .clock(tags_25_clock),
    .reset(tags_25_reset)
  );
  FF_558 tags_26 (
    .clock(tags_26_clock),
    .reset(tags_26_reset)
  );
  FF_558 tags_27 (
    .clock(tags_27_clock),
    .reset(tags_27_reset)
  );
  FF_558 tags_28 (
    .clock(tags_28_clock),
    .reset(tags_28_reset)
  );
  FF_558 tags_29 (
    .clock(tags_29_clock),
    .reset(tags_29_reset)
  );
  FF_558 tags_30 (
    .clock(tags_30_clock),
    .reset(tags_30_reset)
  );
  FF_558 tags_31 (
    .clock(tags_31_clock),
    .reset(tags_31_reset)
  );
  FF_558 tags_32 (
    .clock(tags_32_clock),
    .reset(tags_32_reset)
  );
  FF_558 tags_33 (
    .clock(tags_33_clock),
    .reset(tags_33_reset)
  );
  FF_558 tags_34 (
    .clock(tags_34_clock),
    .reset(tags_34_reset)
  );
  FF_558 tags_35 (
    .clock(tags_35_clock),
    .reset(tags_35_reset)
  );
  FF_558 tags_36 (
    .clock(tags_36_clock),
    .reset(tags_36_reset)
  );
  FF_558 tags_37 (
    .clock(tags_37_clock),
    .reset(tags_37_reset)
  );
  FF_558 tags_38 (
    .clock(tags_38_clock),
    .reset(tags_38_reset)
  );
  FF_558 tags_39 (
    .clock(tags_39_clock),
    .reset(tags_39_reset)
  );
  FF_558 tags_40 (
    .clock(tags_40_clock),
    .reset(tags_40_reset)
  );
  FF_558 tags_41 (
    .clock(tags_41_clock),
    .reset(tags_41_reset)
  );
  FF_558 tags_42 (
    .clock(tags_42_clock),
    .reset(tags_42_reset)
  );
  FF_558 tags_43 (
    .clock(tags_43_clock),
    .reset(tags_43_reset)
  );
  FF_558 tags_44 (
    .clock(tags_44_clock),
    .reset(tags_44_reset)
  );
  FF_558 tags_45 (
    .clock(tags_45_clock),
    .reset(tags_45_reset)
  );
  FF_558 tags_46 (
    .clock(tags_46_clock),
    .reset(tags_46_reset)
  );
  FF_558 tags_47 (
    .clock(tags_47_clock),
    .reset(tags_47_reset)
  );
  FF_558 tags_48 (
    .clock(tags_48_clock),
    .reset(tags_48_reset)
  );
  FF_558 tags_49 (
    .clock(tags_49_clock),
    .reset(tags_49_reset)
  );
  FF_558 tags_50 (
    .clock(tags_50_clock),
    .reset(tags_50_reset)
  );
  FF_558 tags_51 (
    .clock(tags_51_clock),
    .reset(tags_51_reset)
  );
  FF_558 tags_52 (
    .clock(tags_52_clock),
    .reset(tags_52_reset)
  );
  FF_558 tags_53 (
    .clock(tags_53_clock),
    .reset(tags_53_reset)
  );
  FF_558 tags_54 (
    .clock(tags_54_clock),
    .reset(tags_54_reset)
  );
  FF_558 tags_55 (
    .clock(tags_55_clock),
    .reset(tags_55_reset)
  );
  FF_558 tags_56 (
    .clock(tags_56_clock),
    .reset(tags_56_reset)
  );
  FF_558 tags_57 (
    .clock(tags_57_clock),
    .reset(tags_57_reset)
  );
  FF_558 tags_58 (
    .clock(tags_58_clock),
    .reset(tags_58_reset)
  );
  FF_558 tags_59 (
    .clock(tags_59_clock),
    .reset(tags_59_reset)
  );
  FF_558 tags_60 (
    .clock(tags_60_clock),
    .reset(tags_60_reset)
  );
  FF_558 tags_61 (
    .clock(tags_61_clock),
    .reset(tags_61_reset)
  );
  FF_558 tags_62 (
    .clock(tags_62_clock),
    .reset(tags_62_reset)
  );
  FF_558 tags_63 (
    .clock(tags_63_clock),
    .reset(tags_63_reset)
  );
  FF_558 tags_64 (
    .clock(tags_64_clock),
    .reset(tags_64_reset)
  );
  FF_558 tags_65 (
    .clock(tags_65_clock),
    .reset(tags_65_reset)
  );
  FF_558 tags_66 (
    .clock(tags_66_clock),
    .reset(tags_66_reset)
  );
  FF_558 tags_67 (
    .clock(tags_67_clock),
    .reset(tags_67_reset)
  );
  FF_558 tags_68 (
    .clock(tags_68_clock),
    .reset(tags_68_reset)
  );
  FF_558 tags_69 (
    .clock(tags_69_clock),
    .reset(tags_69_reset)
  );
  FF_558 tags_70 (
    .clock(tags_70_clock),
    .reset(tags_70_reset)
  );
  FF_558 tags_71 (
    .clock(tags_71_clock),
    .reset(tags_71_reset)
  );
  FF_558 tags_72 (
    .clock(tags_72_clock),
    .reset(tags_72_reset)
  );
  FF_558 tags_73 (
    .clock(tags_73_clock),
    .reset(tags_73_reset)
  );
  FF_558 tags_74 (
    .clock(tags_74_clock),
    .reset(tags_74_reset)
  );
  FF_558 tags_75 (
    .clock(tags_75_clock),
    .reset(tags_75_reset)
  );
  FF_558 tags_76 (
    .clock(tags_76_clock),
    .reset(tags_76_reset)
  );
  FF_558 tags_77 (
    .clock(tags_77_clock),
    .reset(tags_77_reset)
  );
  FF_558 tags_78 (
    .clock(tags_78_clock),
    .reset(tags_78_reset)
  );
  FF_558 tags_79 (
    .clock(tags_79_clock),
    .reset(tags_79_reset)
  );
  FF_558 tags_80 (
    .clock(tags_80_clock),
    .reset(tags_80_reset)
  );
  FF_558 tags_81 (
    .clock(tags_81_clock),
    .reset(tags_81_reset)
  );
  FF_558 tags_82 (
    .clock(tags_82_clock),
    .reset(tags_82_reset)
  );
  FF_558 tags_83 (
    .clock(tags_83_clock),
    .reset(tags_83_reset)
  );
  FF_558 tags_84 (
    .clock(tags_84_clock),
    .reset(tags_84_reset)
  );
  FF_558 tags_85 (
    .clock(tags_85_clock),
    .reset(tags_85_reset)
  );
  FF_558 tags_86 (
    .clock(tags_86_clock),
    .reset(tags_86_reset)
  );
  FF_558 tags_87 (
    .clock(tags_87_clock),
    .reset(tags_87_reset)
  );
  FF_558 tags_88 (
    .clock(tags_88_clock),
    .reset(tags_88_reset)
  );
  FF_558 tags_89 (
    .clock(tags_89_clock),
    .reset(tags_89_reset)
  );
  FF_558 tags_90 (
    .clock(tags_90_clock),
    .reset(tags_90_reset)
  );
  FF_558 tags_91 (
    .clock(tags_91_clock),
    .reset(tags_91_reset)
  );
  FF_558 tags_92 (
    .clock(tags_92_clock),
    .reset(tags_92_reset)
  );
  FF_558 tags_93 (
    .clock(tags_93_clock),
    .reset(tags_93_reset)
  );
  FF_558 tags_94 (
    .clock(tags_94_clock),
    .reset(tags_94_reset)
  );
  FF_558 tags_95 (
    .clock(tags_95_clock),
    .reset(tags_95_reset)
  );
  FF_558 tags_96 (
    .clock(tags_96_clock),
    .reset(tags_96_reset)
  );
  FF_558 tags_97 (
    .clock(tags_97_clock),
    .reset(tags_97_reset)
  );
  FF_558 tags_98 (
    .clock(tags_98_clock),
    .reset(tags_98_reset)
  );
  FF_558 tags_99 (
    .clock(tags_99_clock),
    .reset(tags_99_reset)
  );
  FF_558 tags_100 (
    .clock(tags_100_clock),
    .reset(tags_100_reset)
  );
  FF_558 tags_101 (
    .clock(tags_101_clock),
    .reset(tags_101_reset)
  );
  FF_558 tags_102 (
    .clock(tags_102_clock),
    .reset(tags_102_reset)
  );
  FF_558 tags_103 (
    .clock(tags_103_clock),
    .reset(tags_103_reset)
  );
  FF_558 tags_104 (
    .clock(tags_104_clock),
    .reset(tags_104_reset)
  );
  FF_558 tags_105 (
    .clock(tags_105_clock),
    .reset(tags_105_reset)
  );
  FF_558 tags_106 (
    .clock(tags_106_clock),
    .reset(tags_106_reset)
  );
  FF_558 tags_107 (
    .clock(tags_107_clock),
    .reset(tags_107_reset)
  );
  FF_558 tags_108 (
    .clock(tags_108_clock),
    .reset(tags_108_reset)
  );
  FF_558 tags_109 (
    .clock(tags_109_clock),
    .reset(tags_109_reset)
  );
  FF_558 tags_110 (
    .clock(tags_110_clock),
    .reset(tags_110_reset)
  );
  FF_558 tags_111 (
    .clock(tags_111_clock),
    .reset(tags_111_reset)
  );
  FF_558 tags_112 (
    .clock(tags_112_clock),
    .reset(tags_112_reset)
  );
  FF_558 tags_113 (
    .clock(tags_113_clock),
    .reset(tags_113_reset)
  );
  FF_558 tags_114 (
    .clock(tags_114_clock),
    .reset(tags_114_reset)
  );
  FF_558 tags_115 (
    .clock(tags_115_clock),
    .reset(tags_115_reset)
  );
  FF_558 tags_116 (
    .clock(tags_116_clock),
    .reset(tags_116_reset)
  );
  FF_558 tags_117 (
    .clock(tags_117_clock),
    .reset(tags_117_reset)
  );
  FF_558 tags_118 (
    .clock(tags_118_clock),
    .reset(tags_118_reset)
  );
  FF_558 tags_119 (
    .clock(tags_119_clock),
    .reset(tags_119_reset)
  );
  FF_558 tags_120 (
    .clock(tags_120_clock),
    .reset(tags_120_reset)
  );
  FF_558 tags_121 (
    .clock(tags_121_clock),
    .reset(tags_121_reset)
  );
  FF_558 tags_122 (
    .clock(tags_122_clock),
    .reset(tags_122_reset)
  );
  FF_558 tags_123 (
    .clock(tags_123_clock),
    .reset(tags_123_reset)
  );
  FF_558 tags_124 (
    .clock(tags_124_clock),
    .reset(tags_124_reset)
  );
  FF_558 tags_125 (
    .clock(tags_125_clock),
    .reset(tags_125_reset)
  );
  FF_558 tags_126 (
    .clock(tags_126_clock),
    .reset(tags_126_reset)
  );
  FF_558 tags_127 (
    .clock(tags_127_clock),
    .reset(tags_127_reset)
  );
  FF_558 tags_128 (
    .clock(tags_128_clock),
    .reset(tags_128_reset)
  );
  FF_558 tags_129 (
    .clock(tags_129_clock),
    .reset(tags_129_reset)
  );
  FF_558 tags_130 (
    .clock(tags_130_clock),
    .reset(tags_130_reset)
  );
  FF_558 tags_131 (
    .clock(tags_131_clock),
    .reset(tags_131_reset)
  );
  FF_558 tags_132 (
    .clock(tags_132_clock),
    .reset(tags_132_reset)
  );
  FF_558 tags_133 (
    .clock(tags_133_clock),
    .reset(tags_133_reset)
  );
  FF_558 tags_134 (
    .clock(tags_134_clock),
    .reset(tags_134_reset)
  );
  FF_558 tags_135 (
    .clock(tags_135_clock),
    .reset(tags_135_reset)
  );
  FF_558 tags_136 (
    .clock(tags_136_clock),
    .reset(tags_136_reset)
  );
  FF_558 tags_137 (
    .clock(tags_137_clock),
    .reset(tags_137_reset)
  );
  FF_558 tags_138 (
    .clock(tags_138_clock),
    .reset(tags_138_reset)
  );
  FF_558 tags_139 (
    .clock(tags_139_clock),
    .reset(tags_139_reset)
  );
  FF_558 tags_140 (
    .clock(tags_140_clock),
    .reset(tags_140_reset)
  );
  FF_558 tags_141 (
    .clock(tags_141_clock),
    .reset(tags_141_reset)
  );
  FF_558 tags_142 (
    .clock(tags_142_clock),
    .reset(tags_142_reset)
  );
  FF_558 tags_143 (
    .clock(tags_143_clock),
    .reset(tags_143_reset)
  );
  FF_558 tags_144 (
    .clock(tags_144_clock),
    .reset(tags_144_reset)
  );
  FF_558 tags_145 (
    .clock(tags_145_clock),
    .reset(tags_145_reset)
  );
  FF_558 tags_146 (
    .clock(tags_146_clock),
    .reset(tags_146_reset)
  );
  FF_558 tags_147 (
    .clock(tags_147_clock),
    .reset(tags_147_reset)
  );
  FF_558 tags_148 (
    .clock(tags_148_clock),
    .reset(tags_148_reset)
  );
  FF_558 tags_149 (
    .clock(tags_149_clock),
    .reset(tags_149_reset)
  );
  FF_558 tags_150 (
    .clock(tags_150_clock),
    .reset(tags_150_reset)
  );
  FF_558 tags_151 (
    .clock(tags_151_clock),
    .reset(tags_151_reset)
  );
  FF_558 tags_152 (
    .clock(tags_152_clock),
    .reset(tags_152_reset)
  );
  FF_558 tags_153 (
    .clock(tags_153_clock),
    .reset(tags_153_reset)
  );
  FF_558 tags_154 (
    .clock(tags_154_clock),
    .reset(tags_154_reset)
  );
  FF_558 tags_155 (
    .clock(tags_155_clock),
    .reset(tags_155_reset)
  );
  FF_558 tags_156 (
    .clock(tags_156_clock),
    .reset(tags_156_reset)
  );
  FF_558 tags_157 (
    .clock(tags_157_clock),
    .reset(tags_157_reset)
  );
  FF_558 tags_158 (
    .clock(tags_158_clock),
    .reset(tags_158_reset)
  );
  FF_558 tags_159 (
    .clock(tags_159_clock),
    .reset(tags_159_reset)
  );
  FF_558 tags_160 (
    .clock(tags_160_clock),
    .reset(tags_160_reset)
  );
  FF_558 tags_161 (
    .clock(tags_161_clock),
    .reset(tags_161_reset)
  );
  FF_558 tags_162 (
    .clock(tags_162_clock),
    .reset(tags_162_reset)
  );
  FF_558 tags_163 (
    .clock(tags_163_clock),
    .reset(tags_163_reset)
  );
  FF_558 tags_164 (
    .clock(tags_164_clock),
    .reset(tags_164_reset)
  );
  FF_558 tags_165 (
    .clock(tags_165_clock),
    .reset(tags_165_reset)
  );
  FF_558 tags_166 (
    .clock(tags_166_clock),
    .reset(tags_166_reset)
  );
  FF_558 tags_167 (
    .clock(tags_167_clock),
    .reset(tags_167_reset)
  );
  FF_558 tags_168 (
    .clock(tags_168_clock),
    .reset(tags_168_reset)
  );
  FF_558 tags_169 (
    .clock(tags_169_clock),
    .reset(tags_169_reset)
  );
  FF_558 tags_170 (
    .clock(tags_170_clock),
    .reset(tags_170_reset)
  );
  FF_558 tags_171 (
    .clock(tags_171_clock),
    .reset(tags_171_reset)
  );
  FF_558 tags_172 (
    .clock(tags_172_clock),
    .reset(tags_172_reset)
  );
  FF_558 tags_173 (
    .clock(tags_173_clock),
    .reset(tags_173_reset)
  );
  FF_558 tags_174 (
    .clock(tags_174_clock),
    .reset(tags_174_reset)
  );
  FF_558 tags_175 (
    .clock(tags_175_clock),
    .reset(tags_175_reset)
  );
  FF_558 tags_176 (
    .clock(tags_176_clock),
    .reset(tags_176_reset)
  );
  FF_558 tags_177 (
    .clock(tags_177_clock),
    .reset(tags_177_reset)
  );
  FF_558 tags_178 (
    .clock(tags_178_clock),
    .reset(tags_178_reset)
  );
  FF_558 tags_179 (
    .clock(tags_179_clock),
    .reset(tags_179_reset)
  );
  FF_558 tags_180 (
    .clock(tags_180_clock),
    .reset(tags_180_reset)
  );
  FF_558 tags_181 (
    .clock(tags_181_clock),
    .reset(tags_181_reset)
  );
  FF_558 tags_182 (
    .clock(tags_182_clock),
    .reset(tags_182_reset)
  );
  FF_558 tags_183 (
    .clock(tags_183_clock),
    .reset(tags_183_reset)
  );
  FF_558 tags_184 (
    .clock(tags_184_clock),
    .reset(tags_184_reset)
  );
  FF_558 tags_185 (
    .clock(tags_185_clock),
    .reset(tags_185_reset)
  );
  FF_558 tags_186 (
    .clock(tags_186_clock),
    .reset(tags_186_reset)
  );
  FF_558 tags_187 (
    .clock(tags_187_clock),
    .reset(tags_187_reset)
  );
  FF_558 tags_188 (
    .clock(tags_188_clock),
    .reset(tags_188_reset)
  );
  FF_558 tags_189 (
    .clock(tags_189_clock),
    .reset(tags_189_reset)
  );
  FF_558 tags_190 (
    .clock(tags_190_clock),
    .reset(tags_190_reset)
  );
  FF_558 tags_191 (
    .clock(tags_191_clock),
    .reset(tags_191_reset)
  );
  FF_558 tags_192 (
    .clock(tags_192_clock),
    .reset(tags_192_reset)
  );
  FF_558 tags_193 (
    .clock(tags_193_clock),
    .reset(tags_193_reset)
  );
  FF_558 tags_194 (
    .clock(tags_194_clock),
    .reset(tags_194_reset)
  );
  FF_558 tags_195 (
    .clock(tags_195_clock),
    .reset(tags_195_reset)
  );
  FF_558 tags_196 (
    .clock(tags_196_clock),
    .reset(tags_196_reset)
  );
  FF_558 tags_197 (
    .clock(tags_197_clock),
    .reset(tags_197_reset)
  );
  FF_558 tags_198 (
    .clock(tags_198_clock),
    .reset(tags_198_reset)
  );
  FF_558 tags_199 (
    .clock(tags_199_clock),
    .reset(tags_199_reset)
  );
  FF_558 tags_200 (
    .clock(tags_200_clock),
    .reset(tags_200_reset)
  );
  FF_558 tags_201 (
    .clock(tags_201_clock),
    .reset(tags_201_reset)
  );
  FF_558 tags_202 (
    .clock(tags_202_clock),
    .reset(tags_202_reset)
  );
  FF_558 tags_203 (
    .clock(tags_203_clock),
    .reset(tags_203_reset)
  );
  FF_558 tags_204 (
    .clock(tags_204_clock),
    .reset(tags_204_reset)
  );
  FF_558 tags_205 (
    .clock(tags_205_clock),
    .reset(tags_205_reset)
  );
  FF_558 tags_206 (
    .clock(tags_206_clock),
    .reset(tags_206_reset)
  );
  FF_558 tags_207 (
    .clock(tags_207_clock),
    .reset(tags_207_reset)
  );
  FF_558 tags_208 (
    .clock(tags_208_clock),
    .reset(tags_208_reset)
  );
  FF_558 tags_209 (
    .clock(tags_209_clock),
    .reset(tags_209_reset)
  );
  FF_558 tags_210 (
    .clock(tags_210_clock),
    .reset(tags_210_reset)
  );
  FF_558 tags_211 (
    .clock(tags_211_clock),
    .reset(tags_211_reset)
  );
  FF_558 tags_212 (
    .clock(tags_212_clock),
    .reset(tags_212_reset)
  );
  FF_558 tags_213 (
    .clock(tags_213_clock),
    .reset(tags_213_reset)
  );
  FF_558 tags_214 (
    .clock(tags_214_clock),
    .reset(tags_214_reset)
  );
  FF_558 tags_215 (
    .clock(tags_215_clock),
    .reset(tags_215_reset)
  );
  FF_558 tags_216 (
    .clock(tags_216_clock),
    .reset(tags_216_reset)
  );
  FF_558 tags_217 (
    .clock(tags_217_clock),
    .reset(tags_217_reset)
  );
  FF_558 tags_218 (
    .clock(tags_218_clock),
    .reset(tags_218_reset)
  );
  FF_558 tags_219 (
    .clock(tags_219_clock),
    .reset(tags_219_reset)
  );
  FF_558 tags_220 (
    .clock(tags_220_clock),
    .reset(tags_220_reset)
  );
  FF_558 tags_221 (
    .clock(tags_221_clock),
    .reset(tags_221_reset)
  );
  FF_558 tags_222 (
    .clock(tags_222_clock),
    .reset(tags_222_reset)
  );
  FF_558 tags_223 (
    .clock(tags_223_clock),
    .reset(tags_223_reset)
  );
  FF_558 tags_224 (
    .clock(tags_224_clock),
    .reset(tags_224_reset)
  );
  FF_558 tags_225 (
    .clock(tags_225_clock),
    .reset(tags_225_reset)
  );
  FF_558 tags_226 (
    .clock(tags_226_clock),
    .reset(tags_226_reset)
  );
  FF_558 tags_227 (
    .clock(tags_227_clock),
    .reset(tags_227_reset)
  );
  FF_558 tags_228 (
    .clock(tags_228_clock),
    .reset(tags_228_reset)
  );
  FF_558 tags_229 (
    .clock(tags_229_clock),
    .reset(tags_229_reset)
  );
  FF_558 tags_230 (
    .clock(tags_230_clock),
    .reset(tags_230_reset)
  );
  FF_558 tags_231 (
    .clock(tags_231_clock),
    .reset(tags_231_reset)
  );
  FF_558 tags_232 (
    .clock(tags_232_clock),
    .reset(tags_232_reset)
  );
  FF_558 tags_233 (
    .clock(tags_233_clock),
    .reset(tags_233_reset)
  );
  FF_558 tags_234 (
    .clock(tags_234_clock),
    .reset(tags_234_reset)
  );
  FF_558 tags_235 (
    .clock(tags_235_clock),
    .reset(tags_235_reset)
  );
  FF_558 tags_236 (
    .clock(tags_236_clock),
    .reset(tags_236_reset)
  );
  FF_558 tags_237 (
    .clock(tags_237_clock),
    .reset(tags_237_reset)
  );
  FF_558 tags_238 (
    .clock(tags_238_clock),
    .reset(tags_238_reset)
  );
  FF_558 tags_239 (
    .clock(tags_239_clock),
    .reset(tags_239_reset)
  );
  FF_558 tags_240 (
    .clock(tags_240_clock),
    .reset(tags_240_reset)
  );
  FF_558 tags_241 (
    .clock(tags_241_clock),
    .reset(tags_241_reset)
  );
  FF_558 tags_242 (
    .clock(tags_242_clock),
    .reset(tags_242_reset)
  );
  FF_558 tags_243 (
    .clock(tags_243_clock),
    .reset(tags_243_reset)
  );
  FF_558 tags_244 (
    .clock(tags_244_clock),
    .reset(tags_244_reset)
  );
  FF_558 tags_245 (
    .clock(tags_245_clock),
    .reset(tags_245_reset)
  );
  FF_558 tags_246 (
    .clock(tags_246_clock),
    .reset(tags_246_reset)
  );
  FF_558 tags_247 (
    .clock(tags_247_clock),
    .reset(tags_247_reset)
  );
  FF_558 tags_248 (
    .clock(tags_248_clock),
    .reset(tags_248_reset)
  );
  FF_558 tags_249 (
    .clock(tags_249_clock),
    .reset(tags_249_reset)
  );
  FF_558 tags_250 (
    .clock(tags_250_clock),
    .reset(tags_250_reset)
  );
  FF_558 tags_251 (
    .clock(tags_251_clock),
    .reset(tags_251_reset)
  );
  FF_558 tags_252 (
    .clock(tags_252_clock),
    .reset(tags_252_reset)
  );
  FF_558 tags_253 (
    .clock(tags_253_clock),
    .reset(tags_253_reset)
  );
  FF_558 tags_254 (
    .clock(tags_254_clock),
    .reset(tags_254_reset)
  );
  FF_558 tags_255 (
    .clock(tags_255_clock),
    .reset(tags_255_reset)
  );
  FF_558 tags_256 (
    .clock(tags_256_clock),
    .reset(tags_256_reset)
  );
  FF_558 tags_257 (
    .clock(tags_257_clock),
    .reset(tags_257_reset)
  );
  FF_558 tags_258 (
    .clock(tags_258_clock),
    .reset(tags_258_reset)
  );
  FF_558 tags_259 (
    .clock(tags_259_clock),
    .reset(tags_259_reset)
  );
  FF_558 tags_260 (
    .clock(tags_260_clock),
    .reset(tags_260_reset)
  );
  FF_558 tags_261 (
    .clock(tags_261_clock),
    .reset(tags_261_reset)
  );
  FF_558 tags_262 (
    .clock(tags_262_clock),
    .reset(tags_262_reset)
  );
  FF_558 tags_263 (
    .clock(tags_263_clock),
    .reset(tags_263_reset)
  );
  FF_558 tags_264 (
    .clock(tags_264_clock),
    .reset(tags_264_reset)
  );
  FF_558 tags_265 (
    .clock(tags_265_clock),
    .reset(tags_265_reset)
  );
  FF_558 tags_266 (
    .clock(tags_266_clock),
    .reset(tags_266_reset)
  );
  FF_558 tags_267 (
    .clock(tags_267_clock),
    .reset(tags_267_reset)
  );
  FF_558 tags_268 (
    .clock(tags_268_clock),
    .reset(tags_268_reset)
  );
  FF_558 tags_269 (
    .clock(tags_269_clock),
    .reset(tags_269_reset)
  );
  FF_558 tags_270 (
    .clock(tags_270_clock),
    .reset(tags_270_reset)
  );
  FF_558 tags_271 (
    .clock(tags_271_clock),
    .reset(tags_271_reset)
  );
  FF_558 tags_272 (
    .clock(tags_272_clock),
    .reset(tags_272_reset)
  );
  FF_558 tags_273 (
    .clock(tags_273_clock),
    .reset(tags_273_reset)
  );
  FF_558 tags_274 (
    .clock(tags_274_clock),
    .reset(tags_274_reset)
  );
  FF_558 tags_275 (
    .clock(tags_275_clock),
    .reset(tags_275_reset)
  );
  FF_558 tags_276 (
    .clock(tags_276_clock),
    .reset(tags_276_reset)
  );
  FF_558 tags_277 (
    .clock(tags_277_clock),
    .reset(tags_277_reset)
  );
  FF_558 tags_278 (
    .clock(tags_278_clock),
    .reset(tags_278_reset)
  );
  FF_558 tags_279 (
    .clock(tags_279_clock),
    .reset(tags_279_reset)
  );
  FF_558 tags_280 (
    .clock(tags_280_clock),
    .reset(tags_280_reset)
  );
  FF_558 tags_281 (
    .clock(tags_281_clock),
    .reset(tags_281_reset)
  );
  FF_558 tags_282 (
    .clock(tags_282_clock),
    .reset(tags_282_reset)
  );
  FF_558 tags_283 (
    .clock(tags_283_clock),
    .reset(tags_283_reset)
  );
  FF_558 tags_284 (
    .clock(tags_284_clock),
    .reset(tags_284_reset)
  );
  FF_558 tags_285 (
    .clock(tags_285_clock),
    .reset(tags_285_reset)
  );
  FF_558 tags_286 (
    .clock(tags_286_clock),
    .reset(tags_286_reset)
  );
  FF_558 tags_287 (
    .clock(tags_287_clock),
    .reset(tags_287_reset)
  );
  FF_558 tags_288 (
    .clock(tags_288_clock),
    .reset(tags_288_reset)
  );
  FF_558 tags_289 (
    .clock(tags_289_clock),
    .reset(tags_289_reset)
  );
  FF_558 tags_290 (
    .clock(tags_290_clock),
    .reset(tags_290_reset)
  );
  FF_558 tags_291 (
    .clock(tags_291_clock),
    .reset(tags_291_reset)
  );
  FF_558 tags_292 (
    .clock(tags_292_clock),
    .reset(tags_292_reset)
  );
  FF_558 tags_293 (
    .clock(tags_293_clock),
    .reset(tags_293_reset)
  );
  FF_558 tags_294 (
    .clock(tags_294_clock),
    .reset(tags_294_reset)
  );
  FF_558 tags_295 (
    .clock(tags_295_clock),
    .reset(tags_295_reset)
  );
  FF_558 tags_296 (
    .clock(tags_296_clock),
    .reset(tags_296_reset)
  );
  FF_558 tags_297 (
    .clock(tags_297_clock),
    .reset(tags_297_reset)
  );
  FF_558 tags_298 (
    .clock(tags_298_clock),
    .reset(tags_298_reset)
  );
  FF_558 tags_299 (
    .clock(tags_299_clock),
    .reset(tags_299_reset)
  );
  FF_558 tags_300 (
    .clock(tags_300_clock),
    .reset(tags_300_reset)
  );
  FF_558 tags_301 (
    .clock(tags_301_clock),
    .reset(tags_301_reset)
  );
  FF_558 tags_302 (
    .clock(tags_302_clock),
    .reset(tags_302_reset)
  );
  FF_558 tags_303 (
    .clock(tags_303_clock),
    .reset(tags_303_reset)
  );
  FF_558 tags_304 (
    .clock(tags_304_clock),
    .reset(tags_304_reset)
  );
  FF_558 tags_305 (
    .clock(tags_305_clock),
    .reset(tags_305_reset)
  );
  FF_558 tags_306 (
    .clock(tags_306_clock),
    .reset(tags_306_reset)
  );
  FF_558 tags_307 (
    .clock(tags_307_clock),
    .reset(tags_307_reset)
  );
  FF_558 tags_308 (
    .clock(tags_308_clock),
    .reset(tags_308_reset)
  );
  FF_558 tags_309 (
    .clock(tags_309_clock),
    .reset(tags_309_reset)
  );
  FF_558 tags_310 (
    .clock(tags_310_clock),
    .reset(tags_310_reset)
  );
  FF_558 tags_311 (
    .clock(tags_311_clock),
    .reset(tags_311_reset)
  );
  FF_558 tags_312 (
    .clock(tags_312_clock),
    .reset(tags_312_reset)
  );
  FF_558 tags_313 (
    .clock(tags_313_clock),
    .reset(tags_313_reset)
  );
  FF_558 tags_314 (
    .clock(tags_314_clock),
    .reset(tags_314_reset)
  );
  FF_558 tags_315 (
    .clock(tags_315_clock),
    .reset(tags_315_reset)
  );
  FF_558 tags_316 (
    .clock(tags_316_clock),
    .reset(tags_316_reset)
  );
  FF_558 tags_317 (
    .clock(tags_317_clock),
    .reset(tags_317_reset)
  );
  FF_558 tags_318 (
    .clock(tags_318_clock),
    .reset(tags_318_reset)
  );
  FF_558 tags_319 (
    .clock(tags_319_clock),
    .reset(tags_319_reset)
  );
  FF_558 tags_320 (
    .clock(tags_320_clock),
    .reset(tags_320_reset)
  );
  FF_558 tags_321 (
    .clock(tags_321_clock),
    .reset(tags_321_reset)
  );
  FF_558 tags_322 (
    .clock(tags_322_clock),
    .reset(tags_322_reset)
  );
  FF_558 tags_323 (
    .clock(tags_323_clock),
    .reset(tags_323_reset)
  );
  FF_558 tags_324 (
    .clock(tags_324_clock),
    .reset(tags_324_reset)
  );
  FF_558 tags_325 (
    .clock(tags_325_clock),
    .reset(tags_325_reset)
  );
  FF_558 tags_326 (
    .clock(tags_326_clock),
    .reset(tags_326_reset)
  );
  FF_558 tags_327 (
    .clock(tags_327_clock),
    .reset(tags_327_reset)
  );
  FF_558 tags_328 (
    .clock(tags_328_clock),
    .reset(tags_328_reset)
  );
  FF_558 tags_329 (
    .clock(tags_329_clock),
    .reset(tags_329_reset)
  );
  FF_558 tags_330 (
    .clock(tags_330_clock),
    .reset(tags_330_reset)
  );
  FF_558 tags_331 (
    .clock(tags_331_clock),
    .reset(tags_331_reset)
  );
  FF_558 tags_332 (
    .clock(tags_332_clock),
    .reset(tags_332_reset)
  );
  FF_558 tags_333 (
    .clock(tags_333_clock),
    .reset(tags_333_reset)
  );
  FF_558 tags_334 (
    .clock(tags_334_clock),
    .reset(tags_334_reset)
  );
  FF_558 tags_335 (
    .clock(tags_335_clock),
    .reset(tags_335_reset)
  );
  FF_558 tags_336 (
    .clock(tags_336_clock),
    .reset(tags_336_reset)
  );
  FF_558 tags_337 (
    .clock(tags_337_clock),
    .reset(tags_337_reset)
  );
  FF_558 tags_338 (
    .clock(tags_338_clock),
    .reset(tags_338_reset)
  );
  FF_558 tags_339 (
    .clock(tags_339_clock),
    .reset(tags_339_reset)
  );
  FF_558 tags_340 (
    .clock(tags_340_clock),
    .reset(tags_340_reset)
  );
  FF_558 tags_341 (
    .clock(tags_341_clock),
    .reset(tags_341_reset)
  );
  FF_558 tags_342 (
    .clock(tags_342_clock),
    .reset(tags_342_reset)
  );
  FF_558 tags_343 (
    .clock(tags_343_clock),
    .reset(tags_343_reset)
  );
  FF_558 tags_344 (
    .clock(tags_344_clock),
    .reset(tags_344_reset)
  );
  FF_558 tags_345 (
    .clock(tags_345_clock),
    .reset(tags_345_reset)
  );
  FF_558 tags_346 (
    .clock(tags_346_clock),
    .reset(tags_346_reset)
  );
  FF_558 tags_347 (
    .clock(tags_347_clock),
    .reset(tags_347_reset)
  );
  FF_558 tags_348 (
    .clock(tags_348_clock),
    .reset(tags_348_reset)
  );
  FF_558 tags_349 (
    .clock(tags_349_clock),
    .reset(tags_349_reset)
  );
  FF_558 tags_350 (
    .clock(tags_350_clock),
    .reset(tags_350_reset)
  );
  FF_558 tags_351 (
    .clock(tags_351_clock),
    .reset(tags_351_reset)
  );
  FF_558 tags_352 (
    .clock(tags_352_clock),
    .reset(tags_352_reset)
  );
  FF_558 tags_353 (
    .clock(tags_353_clock),
    .reset(tags_353_reset)
  );
  FF_558 tags_354 (
    .clock(tags_354_clock),
    .reset(tags_354_reset)
  );
  FF_558 tags_355 (
    .clock(tags_355_clock),
    .reset(tags_355_reset)
  );
  FF_558 tags_356 (
    .clock(tags_356_clock),
    .reset(tags_356_reset)
  );
  FF_558 tags_357 (
    .clock(tags_357_clock),
    .reset(tags_357_reset)
  );
  FF_558 tags_358 (
    .clock(tags_358_clock),
    .reset(tags_358_reset)
  );
  FF_558 tags_359 (
    .clock(tags_359_clock),
    .reset(tags_359_reset)
  );
  FF_558 tags_360 (
    .clock(tags_360_clock),
    .reset(tags_360_reset)
  );
  FF_558 tags_361 (
    .clock(tags_361_clock),
    .reset(tags_361_reset)
  );
  FF_558 tags_362 (
    .clock(tags_362_clock),
    .reset(tags_362_reset)
  );
  FF_558 tags_363 (
    .clock(tags_363_clock),
    .reset(tags_363_reset)
  );
  FF_558 tags_364 (
    .clock(tags_364_clock),
    .reset(tags_364_reset)
  );
  FF_558 tags_365 (
    .clock(tags_365_clock),
    .reset(tags_365_reset)
  );
  FF_558 tags_366 (
    .clock(tags_366_clock),
    .reset(tags_366_reset)
  );
  FF_558 tags_367 (
    .clock(tags_367_clock),
    .reset(tags_367_reset)
  );
  FF_558 tags_368 (
    .clock(tags_368_clock),
    .reset(tags_368_reset)
  );
  FF_558 tags_369 (
    .clock(tags_369_clock),
    .reset(tags_369_reset)
  );
  FF_558 tags_370 (
    .clock(tags_370_clock),
    .reset(tags_370_reset)
  );
  FF_558 tags_371 (
    .clock(tags_371_clock),
    .reset(tags_371_reset)
  );
  FF_558 tags_372 (
    .clock(tags_372_clock),
    .reset(tags_372_reset)
  );
  FF_558 tags_373 (
    .clock(tags_373_clock),
    .reset(tags_373_reset)
  );
  FF_558 tags_374 (
    .clock(tags_374_clock),
    .reset(tags_374_reset)
  );
  FF_558 tags_375 (
    .clock(tags_375_clock),
    .reset(tags_375_reset)
  );
  FF_558 tags_376 (
    .clock(tags_376_clock),
    .reset(tags_376_reset)
  );
  FF_558 tags_377 (
    .clock(tags_377_clock),
    .reset(tags_377_reset)
  );
  FF_558 tags_378 (
    .clock(tags_378_clock),
    .reset(tags_378_reset)
  );
  FF_558 tags_379 (
    .clock(tags_379_clock),
    .reset(tags_379_reset)
  );
  FF_558 tags_380 (
    .clock(tags_380_clock),
    .reset(tags_380_reset)
  );
  FF_558 tags_381 (
    .clock(tags_381_clock),
    .reset(tags_381_reset)
  );
  FF_558 tags_382 (
    .clock(tags_382_clock),
    .reset(tags_382_reset)
  );
  FF_558 tags_383 (
    .clock(tags_383_clock),
    .reset(tags_383_reset)
  );
  FF_558 tags_384 (
    .clock(tags_384_clock),
    .reset(tags_384_reset)
  );
  FF_558 tags_385 (
    .clock(tags_385_clock),
    .reset(tags_385_reset)
  );
  FF_558 tags_386 (
    .clock(tags_386_clock),
    .reset(tags_386_reset)
  );
  FF_558 tags_387 (
    .clock(tags_387_clock),
    .reset(tags_387_reset)
  );
  FF_558 tags_388 (
    .clock(tags_388_clock),
    .reset(tags_388_reset)
  );
  FF_558 tags_389 (
    .clock(tags_389_clock),
    .reset(tags_389_reset)
  );
  FF_558 tags_390 (
    .clock(tags_390_clock),
    .reset(tags_390_reset)
  );
  FF_558 tags_391 (
    .clock(tags_391_clock),
    .reset(tags_391_reset)
  );
  FF_558 tags_392 (
    .clock(tags_392_clock),
    .reset(tags_392_reset)
  );
  FF_558 tags_393 (
    .clock(tags_393_clock),
    .reset(tags_393_reset)
  );
  FF_558 tags_394 (
    .clock(tags_394_clock),
    .reset(tags_394_reset)
  );
  FF_558 tags_395 (
    .clock(tags_395_clock),
    .reset(tags_395_reset)
  );
  FF_558 tags_396 (
    .clock(tags_396_clock),
    .reset(tags_396_reset)
  );
  FF_558 tags_397 (
    .clock(tags_397_clock),
    .reset(tags_397_reset)
  );
  FF_558 tags_398 (
    .clock(tags_398_clock),
    .reset(tags_398_reset)
  );
  FF_558 tags_399 (
    .clock(tags_399_clock),
    .reset(tags_399_reset)
  );
  FF_558 tags_400 (
    .clock(tags_400_clock),
    .reset(tags_400_reset)
  );
  FF_558 tags_401 (
    .clock(tags_401_clock),
    .reset(tags_401_reset)
  );
  FF_558 tags_402 (
    .clock(tags_402_clock),
    .reset(tags_402_reset)
  );
  FF_558 tags_403 (
    .clock(tags_403_clock),
    .reset(tags_403_reset)
  );
  FF_558 tags_404 (
    .clock(tags_404_clock),
    .reset(tags_404_reset)
  );
  FF_558 tags_405 (
    .clock(tags_405_clock),
    .reset(tags_405_reset)
  );
  FF_558 tags_406 (
    .clock(tags_406_clock),
    .reset(tags_406_reset)
  );
  FF_558 tags_407 (
    .clock(tags_407_clock),
    .reset(tags_407_reset)
  );
  FF_558 tags_408 (
    .clock(tags_408_clock),
    .reset(tags_408_reset)
  );
  FF_558 tags_409 (
    .clock(tags_409_clock),
    .reset(tags_409_reset)
  );
  FF_558 tags_410 (
    .clock(tags_410_clock),
    .reset(tags_410_reset)
  );
  FF_558 tags_411 (
    .clock(tags_411_clock),
    .reset(tags_411_reset)
  );
  FF_558 tags_412 (
    .clock(tags_412_clock),
    .reset(tags_412_reset)
  );
  FF_558 tags_413 (
    .clock(tags_413_clock),
    .reset(tags_413_reset)
  );
  FF_558 tags_414 (
    .clock(tags_414_clock),
    .reset(tags_414_reset)
  );
  FF_558 tags_415 (
    .clock(tags_415_clock),
    .reset(tags_415_reset)
  );
  FF_558 tags_416 (
    .clock(tags_416_clock),
    .reset(tags_416_reset)
  );
  FF_558 tags_417 (
    .clock(tags_417_clock),
    .reset(tags_417_reset)
  );
  FF_558 tags_418 (
    .clock(tags_418_clock),
    .reset(tags_418_reset)
  );
  FF_558 tags_419 (
    .clock(tags_419_clock),
    .reset(tags_419_reset)
  );
  FF_558 tags_420 (
    .clock(tags_420_clock),
    .reset(tags_420_reset)
  );
  FF_558 tags_421 (
    .clock(tags_421_clock),
    .reset(tags_421_reset)
  );
  FF_558 tags_422 (
    .clock(tags_422_clock),
    .reset(tags_422_reset)
  );
  FF_558 tags_423 (
    .clock(tags_423_clock),
    .reset(tags_423_reset)
  );
  FF_558 tags_424 (
    .clock(tags_424_clock),
    .reset(tags_424_reset)
  );
  FF_558 tags_425 (
    .clock(tags_425_clock),
    .reset(tags_425_reset)
  );
  FF_558 tags_426 (
    .clock(tags_426_clock),
    .reset(tags_426_reset)
  );
  FF_558 tags_427 (
    .clock(tags_427_clock),
    .reset(tags_427_reset)
  );
  FF_558 tags_428 (
    .clock(tags_428_clock),
    .reset(tags_428_reset)
  );
  FF_558 tags_429 (
    .clock(tags_429_clock),
    .reset(tags_429_reset)
  );
  FF_558 tags_430 (
    .clock(tags_430_clock),
    .reset(tags_430_reset)
  );
  FF_558 tags_431 (
    .clock(tags_431_clock),
    .reset(tags_431_reset)
  );
  FF_558 tags_432 (
    .clock(tags_432_clock),
    .reset(tags_432_reset)
  );
  FF_558 tags_433 (
    .clock(tags_433_clock),
    .reset(tags_433_reset)
  );
  FF_558 tags_434 (
    .clock(tags_434_clock),
    .reset(tags_434_reset)
  );
  FF_558 tags_435 (
    .clock(tags_435_clock),
    .reset(tags_435_reset)
  );
  FF_558 tags_436 (
    .clock(tags_436_clock),
    .reset(tags_436_reset)
  );
  FF_558 tags_437 (
    .clock(tags_437_clock),
    .reset(tags_437_reset)
  );
  FF_558 tags_438 (
    .clock(tags_438_clock),
    .reset(tags_438_reset)
  );
  FF_558 tags_439 (
    .clock(tags_439_clock),
    .reset(tags_439_reset)
  );
  FF_558 tags_440 (
    .clock(tags_440_clock),
    .reset(tags_440_reset)
  );
  FF_558 tags_441 (
    .clock(tags_441_clock),
    .reset(tags_441_reset)
  );
  FF_558 tags_442 (
    .clock(tags_442_clock),
    .reset(tags_442_reset)
  );
  FF_558 tags_443 (
    .clock(tags_443_clock),
    .reset(tags_443_reset)
  );
  FF_558 tags_444 (
    .clock(tags_444_clock),
    .reset(tags_444_reset)
  );
  FF_558 tags_445 (
    .clock(tags_445_clock),
    .reset(tags_445_reset)
  );
  FF_558 tags_446 (
    .clock(tags_446_clock),
    .reset(tags_446_reset)
  );
  FF_558 tags_447 (
    .clock(tags_447_clock),
    .reset(tags_447_reset)
  );
  FF_558 tags_448 (
    .clock(tags_448_clock),
    .reset(tags_448_reset)
  );
  FF_558 tags_449 (
    .clock(tags_449_clock),
    .reset(tags_449_reset)
  );
  FF_558 tags_450 (
    .clock(tags_450_clock),
    .reset(tags_450_reset)
  );
  FF_558 tags_451 (
    .clock(tags_451_clock),
    .reset(tags_451_reset)
  );
  FF_558 tags_452 (
    .clock(tags_452_clock),
    .reset(tags_452_reset)
  );
  FF_558 tags_453 (
    .clock(tags_453_clock),
    .reset(tags_453_reset)
  );
  FF_558 tags_454 (
    .clock(tags_454_clock),
    .reset(tags_454_reset)
  );
  FF_558 tags_455 (
    .clock(tags_455_clock),
    .reset(tags_455_reset)
  );
  FF_558 tags_456 (
    .clock(tags_456_clock),
    .reset(tags_456_reset)
  );
  FF_558 tags_457 (
    .clock(tags_457_clock),
    .reset(tags_457_reset)
  );
  FF_558 tags_458 (
    .clock(tags_458_clock),
    .reset(tags_458_reset)
  );
  FF_558 tags_459 (
    .clock(tags_459_clock),
    .reset(tags_459_reset)
  );
  FF_558 tags_460 (
    .clock(tags_460_clock),
    .reset(tags_460_reset)
  );
  FF_558 tags_461 (
    .clock(tags_461_clock),
    .reset(tags_461_reset)
  );
  FF_558 tags_462 (
    .clock(tags_462_clock),
    .reset(tags_462_reset)
  );
  FF_558 tags_463 (
    .clock(tags_463_clock),
    .reset(tags_463_reset)
  );
  FF_558 tags_464 (
    .clock(tags_464_clock),
    .reset(tags_464_reset)
  );
  FF_558 tags_465 (
    .clock(tags_465_clock),
    .reset(tags_465_reset)
  );
  FF_558 tags_466 (
    .clock(tags_466_clock),
    .reset(tags_466_reset)
  );
  FF_558 tags_467 (
    .clock(tags_467_clock),
    .reset(tags_467_reset)
  );
  FF_558 tags_468 (
    .clock(tags_468_clock),
    .reset(tags_468_reset)
  );
  FF_558 tags_469 (
    .clock(tags_469_clock),
    .reset(tags_469_reset)
  );
  FF_558 tags_470 (
    .clock(tags_470_clock),
    .reset(tags_470_reset)
  );
  FF_558 tags_471 (
    .clock(tags_471_clock),
    .reset(tags_471_reset)
  );
  FF_558 tags_472 (
    .clock(tags_472_clock),
    .reset(tags_472_reset)
  );
  FF_558 tags_473 (
    .clock(tags_473_clock),
    .reset(tags_473_reset)
  );
  FF_558 tags_474 (
    .clock(tags_474_clock),
    .reset(tags_474_reset)
  );
  FF_558 tags_475 (
    .clock(tags_475_clock),
    .reset(tags_475_reset)
  );
  FF_558 tags_476 (
    .clock(tags_476_clock),
    .reset(tags_476_reset)
  );
  FF_558 tags_477 (
    .clock(tags_477_clock),
    .reset(tags_477_reset)
  );
  FF_558 tags_478 (
    .clock(tags_478_clock),
    .reset(tags_478_reset)
  );
  FF_558 tags_479 (
    .clock(tags_479_clock),
    .reset(tags_479_reset)
  );
  FF_558 tags_480 (
    .clock(tags_480_clock),
    .reset(tags_480_reset)
  );
  FF_558 tags_481 (
    .clock(tags_481_clock),
    .reset(tags_481_reset)
  );
  FF_558 tags_482 (
    .clock(tags_482_clock),
    .reset(tags_482_reset)
  );
  FF_558 tags_483 (
    .clock(tags_483_clock),
    .reset(tags_483_reset)
  );
  FF_558 tags_484 (
    .clock(tags_484_clock),
    .reset(tags_484_reset)
  );
  FF_558 tags_485 (
    .clock(tags_485_clock),
    .reset(tags_485_reset)
  );
  FF_558 tags_486 (
    .clock(tags_486_clock),
    .reset(tags_486_reset)
  );
  FF_558 tags_487 (
    .clock(tags_487_clock),
    .reset(tags_487_reset)
  );
  FF_558 tags_488 (
    .clock(tags_488_clock),
    .reset(tags_488_reset)
  );
  FF_558 tags_489 (
    .clock(tags_489_clock),
    .reset(tags_489_reset)
  );
  FF_558 tags_490 (
    .clock(tags_490_clock),
    .reset(tags_490_reset)
  );
  FF_558 tags_491 (
    .clock(tags_491_clock),
    .reset(tags_491_reset)
  );
  FF_558 tags_492 (
    .clock(tags_492_clock),
    .reset(tags_492_reset)
  );
  FF_558 tags_493 (
    .clock(tags_493_clock),
    .reset(tags_493_reset)
  );
  FF_558 tags_494 (
    .clock(tags_494_clock),
    .reset(tags_494_reset)
  );
  FF_558 tags_495 (
    .clock(tags_495_clock),
    .reset(tags_495_reset)
  );
  FF_558 tags_496 (
    .clock(tags_496_clock),
    .reset(tags_496_reset)
  );
  FF_558 tags_497 (
    .clock(tags_497_clock),
    .reset(tags_497_reset)
  );
  FF_558 tags_498 (
    .clock(tags_498_clock),
    .reset(tags_498_reset)
  );
  FF_558 tags_499 (
    .clock(tags_499_clock),
    .reset(tags_499_reset)
  );
  FF_558 tags_500 (
    .clock(tags_500_clock),
    .reset(tags_500_reset)
  );
  FF_558 tags_501 (
    .clock(tags_501_clock),
    .reset(tags_501_reset)
  );
  FF_558 tags_502 (
    .clock(tags_502_clock),
    .reset(tags_502_reset)
  );
  FF_558 tags_503 (
    .clock(tags_503_clock),
    .reset(tags_503_reset)
  );
  FF_558 tags_504 (
    .clock(tags_504_clock),
    .reset(tags_504_reset)
  );
  FF_558 tags_505 (
    .clock(tags_505_clock),
    .reset(tags_505_reset)
  );
  FF_558 tags_506 (
    .clock(tags_506_clock),
    .reset(tags_506_reset)
  );
  FF_558 tags_507 (
    .clock(tags_507_clock),
    .reset(tags_507_reset)
  );
  FF_558 tags_508 (
    .clock(tags_508_clock),
    .reset(tags_508_reset)
  );
  FF_558 tags_509 (
    .clock(tags_509_clock),
    .reset(tags_509_reset)
  );
  FF_558 tags_510 (
    .clock(tags_510_clock),
    .reset(tags_510_reset)
  );
  FF_558 tags_511 (
    .clock(tags_511_clock),
    .reset(tags_511_reset)
  );
  SRAMByteEnable metadata (
    .clock(metadata_clock),
    .io_wdata_0(metadata_io_wdata_0),
    .io_wdata_1(metadata_io_wdata_1),
    .io_wdata_2(metadata_io_wdata_2),
    .io_wdata_3(metadata_io_wdata_3),
    .io_wdata_4(metadata_io_wdata_4),
    .io_wdata_5(metadata_io_wdata_5),
    .io_wdata_6(metadata_io_wdata_6),
    .io_wdata_7(metadata_io_wdata_7),
    .io_wdata_8(metadata_io_wdata_8),
    .io_wdata_9(metadata_io_wdata_9),
    .io_wdata_10(metadata_io_wdata_10),
    .io_wdata_11(metadata_io_wdata_11),
    .io_wdata_12(metadata_io_wdata_12),
    .io_wdata_13(metadata_io_wdata_13),
    .io_wdata_14(metadata_io_wdata_14),
    .io_wdata_15(metadata_io_wdata_15),
    .io_rdata_0(metadata_io_rdata_0),
    .io_rdata_1(metadata_io_rdata_1),
    .io_rdata_2(metadata_io_rdata_2),
    .io_rdata_3(metadata_io_rdata_3),
    .io_rdata_4(metadata_io_rdata_4),
    .io_rdata_5(metadata_io_rdata_5),
    .io_rdata_6(metadata_io_rdata_6),
    .io_rdata_7(metadata_io_rdata_7),
    .io_rdata_8(metadata_io_rdata_8),
    .io_rdata_9(metadata_io_rdata_9),
    .io_rdata_10(metadata_io_rdata_10),
    .io_rdata_11(metadata_io_rdata_11),
    .io_rdata_12(metadata_io_rdata_12),
    .io_rdata_13(metadata_io_rdata_13),
    .io_rdata_14(metadata_io_rdata_14),
    .io_rdata_15(metadata_io_rdata_15)
  );
  assign _T_19089 = io_waddr[5:2];
  assign _T_19127 = {1'h1,woffset};
  assign _GEN_2 = 4'h0 == io_position ? _GEN_0 : 8'h0;
  assign _GEN_3 = 4'h1 == io_position ? _GEN_0 : 8'h0;
  assign _GEN_4 = 4'h2 == io_position ? _GEN_0 : 8'h0;
  assign _GEN_5 = 4'h3 == io_position ? _GEN_0 : 8'h0;
  assign _GEN_6 = 4'h4 == io_position ? _GEN_0 : 8'h0;
  assign _GEN_7 = 4'h5 == io_position ? _GEN_0 : 8'h0;
  assign _GEN_8 = 4'h6 == io_position ? _GEN_0 : 8'h0;
  assign _GEN_9 = 4'h7 == io_position ? _GEN_0 : 8'h0;
  assign _GEN_10 = 4'h8 == io_position ? _GEN_0 : 8'h0;
  assign _GEN_11 = 4'h9 == io_position ? _GEN_0 : 8'h0;
  assign _GEN_12 = 4'ha == io_position ? _GEN_0 : 8'h0;
  assign _GEN_13 = 4'hb == io_position ? _GEN_0 : 8'h0;
  assign _GEN_14 = 4'hc == io_position ? _GEN_0 : 8'h0;
  assign _GEN_15 = 4'hd == io_position ? _GEN_0 : 8'h0;
  assign _GEN_16 = 4'he == io_position ? _GEN_0 : 8'h0;
  assign _GEN_17 = 4'hf == io_position ? _GEN_0 : 8'h0;
  assign io_rmetaData_0 = metadata_io_rdata_0;
  assign io_rmetaData_1 = metadata_io_rdata_1;
  assign io_rmetaData_2 = metadata_io_rdata_2;
  assign io_rmetaData_3 = metadata_io_rdata_3;
  assign io_rmetaData_4 = metadata_io_rdata_4;
  assign io_rmetaData_5 = metadata_io_rdata_5;
  assign io_rmetaData_6 = metadata_io_rdata_6;
  assign io_rmetaData_7 = metadata_io_rdata_7;
  assign io_rmetaData_8 = metadata_io_rdata_8;
  assign io_rmetaData_9 = metadata_io_rdata_9;
  assign io_rmetaData_10 = metadata_io_rdata_10;
  assign io_rmetaData_11 = metadata_io_rdata_11;
  assign io_rmetaData_12 = metadata_io_rdata_12;
  assign io_rmetaData_13 = metadata_io_rdata_13;
  assign io_rmetaData_14 = metadata_io_rdata_14;
  assign io_rmetaData_15 = metadata_io_rdata_15;
  assign valid_0_io_in = 1'h1;
  assign valid_0_io_enable = 1'h0;
  assign valid_0_clock = clock;
  assign valid_0_reset = reset;
  assign valid_1_io_in = 1'h1;
  assign valid_1_io_enable = 1'h0;
  assign valid_1_clock = clock;
  assign valid_1_reset = reset;
  assign valid_2_io_in = 1'h1;
  assign valid_2_io_enable = 1'h0;
  assign valid_2_clock = clock;
  assign valid_2_reset = reset;
  assign valid_3_io_in = 1'h1;
  assign valid_3_io_enable = 1'h0;
  assign valid_3_clock = clock;
  assign valid_3_reset = reset;
  assign valid_4_io_in = 1'h1;
  assign valid_4_io_enable = 1'h0;
  assign valid_4_clock = clock;
  assign valid_4_reset = reset;
  assign valid_5_io_in = 1'h1;
  assign valid_5_io_enable = 1'h0;
  assign valid_5_clock = clock;
  assign valid_5_reset = reset;
  assign valid_6_io_in = 1'h1;
  assign valid_6_io_enable = 1'h0;
  assign valid_6_clock = clock;
  assign valid_6_reset = reset;
  assign valid_7_io_in = 1'h1;
  assign valid_7_io_enable = 1'h0;
  assign valid_7_clock = clock;
  assign valid_7_reset = reset;
  assign valid_8_io_in = 1'h1;
  assign valid_8_io_enable = 1'h0;
  assign valid_8_clock = clock;
  assign valid_8_reset = reset;
  assign valid_9_io_in = 1'h1;
  assign valid_9_io_enable = 1'h0;
  assign valid_9_clock = clock;
  assign valid_9_reset = reset;
  assign valid_10_io_in = 1'h1;
  assign valid_10_io_enable = 1'h0;
  assign valid_10_clock = clock;
  assign valid_10_reset = reset;
  assign valid_11_io_in = 1'h1;
  assign valid_11_io_enable = 1'h0;
  assign valid_11_clock = clock;
  assign valid_11_reset = reset;
  assign valid_12_io_in = 1'h1;
  assign valid_12_io_enable = 1'h0;
  assign valid_12_clock = clock;
  assign valid_12_reset = reset;
  assign valid_13_io_in = 1'h1;
  assign valid_13_io_enable = 1'h0;
  assign valid_13_clock = clock;
  assign valid_13_reset = reset;
  assign valid_14_io_in = 1'h1;
  assign valid_14_io_enable = 1'h0;
  assign valid_14_clock = clock;
  assign valid_14_reset = reset;
  assign valid_15_io_in = 1'h1;
  assign valid_15_io_enable = 1'h0;
  assign valid_15_clock = clock;
  assign valid_15_reset = reset;
  assign valid_16_io_in = 1'h1;
  assign valid_16_io_enable = 1'h0;
  assign valid_16_clock = clock;
  assign valid_16_reset = reset;
  assign valid_17_io_in = 1'h1;
  assign valid_17_io_enable = 1'h0;
  assign valid_17_clock = clock;
  assign valid_17_reset = reset;
  assign valid_18_io_in = 1'h1;
  assign valid_18_io_enable = 1'h0;
  assign valid_18_clock = clock;
  assign valid_18_reset = reset;
  assign valid_19_io_in = 1'h1;
  assign valid_19_io_enable = 1'h0;
  assign valid_19_clock = clock;
  assign valid_19_reset = reset;
  assign valid_20_io_in = 1'h1;
  assign valid_20_io_enable = 1'h0;
  assign valid_20_clock = clock;
  assign valid_20_reset = reset;
  assign valid_21_io_in = 1'h1;
  assign valid_21_io_enable = 1'h0;
  assign valid_21_clock = clock;
  assign valid_21_reset = reset;
  assign valid_22_io_in = 1'h1;
  assign valid_22_io_enable = 1'h0;
  assign valid_22_clock = clock;
  assign valid_22_reset = reset;
  assign valid_23_io_in = 1'h1;
  assign valid_23_io_enable = 1'h0;
  assign valid_23_clock = clock;
  assign valid_23_reset = reset;
  assign valid_24_io_in = 1'h1;
  assign valid_24_io_enable = 1'h0;
  assign valid_24_clock = clock;
  assign valid_24_reset = reset;
  assign valid_25_io_in = 1'h1;
  assign valid_25_io_enable = 1'h0;
  assign valid_25_clock = clock;
  assign valid_25_reset = reset;
  assign valid_26_io_in = 1'h1;
  assign valid_26_io_enable = 1'h0;
  assign valid_26_clock = clock;
  assign valid_26_reset = reset;
  assign valid_27_io_in = 1'h1;
  assign valid_27_io_enable = 1'h0;
  assign valid_27_clock = clock;
  assign valid_27_reset = reset;
  assign valid_28_io_in = 1'h1;
  assign valid_28_io_enable = 1'h0;
  assign valid_28_clock = clock;
  assign valid_28_reset = reset;
  assign valid_29_io_in = 1'h1;
  assign valid_29_io_enable = 1'h0;
  assign valid_29_clock = clock;
  assign valid_29_reset = reset;
  assign valid_30_io_in = 1'h1;
  assign valid_30_io_enable = 1'h0;
  assign valid_30_clock = clock;
  assign valid_30_reset = reset;
  assign valid_31_io_in = 1'h1;
  assign valid_31_io_enable = 1'h0;
  assign valid_31_clock = clock;
  assign valid_31_reset = reset;
  assign valid_32_io_in = 1'h1;
  assign valid_32_io_enable = 1'h0;
  assign valid_32_clock = clock;
  assign valid_32_reset = reset;
  assign valid_33_io_in = 1'h1;
  assign valid_33_io_enable = 1'h0;
  assign valid_33_clock = clock;
  assign valid_33_reset = reset;
  assign valid_34_io_in = 1'h1;
  assign valid_34_io_enable = 1'h0;
  assign valid_34_clock = clock;
  assign valid_34_reset = reset;
  assign valid_35_io_in = 1'h1;
  assign valid_35_io_enable = 1'h0;
  assign valid_35_clock = clock;
  assign valid_35_reset = reset;
  assign valid_36_io_in = 1'h1;
  assign valid_36_io_enable = 1'h0;
  assign valid_36_clock = clock;
  assign valid_36_reset = reset;
  assign valid_37_io_in = 1'h1;
  assign valid_37_io_enable = 1'h0;
  assign valid_37_clock = clock;
  assign valid_37_reset = reset;
  assign valid_38_io_in = 1'h1;
  assign valid_38_io_enable = 1'h0;
  assign valid_38_clock = clock;
  assign valid_38_reset = reset;
  assign valid_39_io_in = 1'h1;
  assign valid_39_io_enable = 1'h0;
  assign valid_39_clock = clock;
  assign valid_39_reset = reset;
  assign valid_40_io_in = 1'h1;
  assign valid_40_io_enable = 1'h0;
  assign valid_40_clock = clock;
  assign valid_40_reset = reset;
  assign valid_41_io_in = 1'h1;
  assign valid_41_io_enable = 1'h0;
  assign valid_41_clock = clock;
  assign valid_41_reset = reset;
  assign valid_42_io_in = 1'h1;
  assign valid_42_io_enable = 1'h0;
  assign valid_42_clock = clock;
  assign valid_42_reset = reset;
  assign valid_43_io_in = 1'h1;
  assign valid_43_io_enable = 1'h0;
  assign valid_43_clock = clock;
  assign valid_43_reset = reset;
  assign valid_44_io_in = 1'h1;
  assign valid_44_io_enable = 1'h0;
  assign valid_44_clock = clock;
  assign valid_44_reset = reset;
  assign valid_45_io_in = 1'h1;
  assign valid_45_io_enable = 1'h0;
  assign valid_45_clock = clock;
  assign valid_45_reset = reset;
  assign valid_46_io_in = 1'h1;
  assign valid_46_io_enable = 1'h0;
  assign valid_46_clock = clock;
  assign valid_46_reset = reset;
  assign valid_47_io_in = 1'h1;
  assign valid_47_io_enable = 1'h0;
  assign valid_47_clock = clock;
  assign valid_47_reset = reset;
  assign valid_48_io_in = 1'h1;
  assign valid_48_io_enable = 1'h0;
  assign valid_48_clock = clock;
  assign valid_48_reset = reset;
  assign valid_49_io_in = 1'h1;
  assign valid_49_io_enable = 1'h0;
  assign valid_49_clock = clock;
  assign valid_49_reset = reset;
  assign valid_50_io_in = 1'h1;
  assign valid_50_io_enable = 1'h0;
  assign valid_50_clock = clock;
  assign valid_50_reset = reset;
  assign valid_51_io_in = 1'h1;
  assign valid_51_io_enable = 1'h0;
  assign valid_51_clock = clock;
  assign valid_51_reset = reset;
  assign valid_52_io_in = 1'h1;
  assign valid_52_io_enable = 1'h0;
  assign valid_52_clock = clock;
  assign valid_52_reset = reset;
  assign valid_53_io_in = 1'h1;
  assign valid_53_io_enable = 1'h0;
  assign valid_53_clock = clock;
  assign valid_53_reset = reset;
  assign valid_54_io_in = 1'h1;
  assign valid_54_io_enable = 1'h0;
  assign valid_54_clock = clock;
  assign valid_54_reset = reset;
  assign valid_55_io_in = 1'h1;
  assign valid_55_io_enable = 1'h0;
  assign valid_55_clock = clock;
  assign valid_55_reset = reset;
  assign valid_56_io_in = 1'h1;
  assign valid_56_io_enable = 1'h0;
  assign valid_56_clock = clock;
  assign valid_56_reset = reset;
  assign valid_57_io_in = 1'h1;
  assign valid_57_io_enable = 1'h0;
  assign valid_57_clock = clock;
  assign valid_57_reset = reset;
  assign valid_58_io_in = 1'h1;
  assign valid_58_io_enable = 1'h0;
  assign valid_58_clock = clock;
  assign valid_58_reset = reset;
  assign valid_59_io_in = 1'h1;
  assign valid_59_io_enable = 1'h0;
  assign valid_59_clock = clock;
  assign valid_59_reset = reset;
  assign valid_60_io_in = 1'h1;
  assign valid_60_io_enable = 1'h0;
  assign valid_60_clock = clock;
  assign valid_60_reset = reset;
  assign valid_61_io_in = 1'h1;
  assign valid_61_io_enable = 1'h0;
  assign valid_61_clock = clock;
  assign valid_61_reset = reset;
  assign valid_62_io_in = 1'h1;
  assign valid_62_io_enable = 1'h0;
  assign valid_62_clock = clock;
  assign valid_62_reset = reset;
  assign valid_63_io_in = 1'h1;
  assign valid_63_io_enable = 1'h0;
  assign valid_63_clock = clock;
  assign valid_63_reset = reset;
  assign valid_64_io_in = 1'h1;
  assign valid_64_io_enable = 1'h0;
  assign valid_64_clock = clock;
  assign valid_64_reset = reset;
  assign valid_65_io_in = 1'h1;
  assign valid_65_io_enable = 1'h0;
  assign valid_65_clock = clock;
  assign valid_65_reset = reset;
  assign valid_66_io_in = 1'h1;
  assign valid_66_io_enable = 1'h0;
  assign valid_66_clock = clock;
  assign valid_66_reset = reset;
  assign valid_67_io_in = 1'h1;
  assign valid_67_io_enable = 1'h0;
  assign valid_67_clock = clock;
  assign valid_67_reset = reset;
  assign valid_68_io_in = 1'h1;
  assign valid_68_io_enable = 1'h0;
  assign valid_68_clock = clock;
  assign valid_68_reset = reset;
  assign valid_69_io_in = 1'h1;
  assign valid_69_io_enable = 1'h0;
  assign valid_69_clock = clock;
  assign valid_69_reset = reset;
  assign valid_70_io_in = 1'h1;
  assign valid_70_io_enable = 1'h0;
  assign valid_70_clock = clock;
  assign valid_70_reset = reset;
  assign valid_71_io_in = 1'h1;
  assign valid_71_io_enable = 1'h0;
  assign valid_71_clock = clock;
  assign valid_71_reset = reset;
  assign valid_72_io_in = 1'h1;
  assign valid_72_io_enable = 1'h0;
  assign valid_72_clock = clock;
  assign valid_72_reset = reset;
  assign valid_73_io_in = 1'h1;
  assign valid_73_io_enable = 1'h0;
  assign valid_73_clock = clock;
  assign valid_73_reset = reset;
  assign valid_74_io_in = 1'h1;
  assign valid_74_io_enable = 1'h0;
  assign valid_74_clock = clock;
  assign valid_74_reset = reset;
  assign valid_75_io_in = 1'h1;
  assign valid_75_io_enable = 1'h0;
  assign valid_75_clock = clock;
  assign valid_75_reset = reset;
  assign valid_76_io_in = 1'h1;
  assign valid_76_io_enable = 1'h0;
  assign valid_76_clock = clock;
  assign valid_76_reset = reset;
  assign valid_77_io_in = 1'h1;
  assign valid_77_io_enable = 1'h0;
  assign valid_77_clock = clock;
  assign valid_77_reset = reset;
  assign valid_78_io_in = 1'h1;
  assign valid_78_io_enable = 1'h0;
  assign valid_78_clock = clock;
  assign valid_78_reset = reset;
  assign valid_79_io_in = 1'h1;
  assign valid_79_io_enable = 1'h0;
  assign valid_79_clock = clock;
  assign valid_79_reset = reset;
  assign valid_80_io_in = 1'h1;
  assign valid_80_io_enable = 1'h0;
  assign valid_80_clock = clock;
  assign valid_80_reset = reset;
  assign valid_81_io_in = 1'h1;
  assign valid_81_io_enable = 1'h0;
  assign valid_81_clock = clock;
  assign valid_81_reset = reset;
  assign valid_82_io_in = 1'h1;
  assign valid_82_io_enable = 1'h0;
  assign valid_82_clock = clock;
  assign valid_82_reset = reset;
  assign valid_83_io_in = 1'h1;
  assign valid_83_io_enable = 1'h0;
  assign valid_83_clock = clock;
  assign valid_83_reset = reset;
  assign valid_84_io_in = 1'h1;
  assign valid_84_io_enable = 1'h0;
  assign valid_84_clock = clock;
  assign valid_84_reset = reset;
  assign valid_85_io_in = 1'h1;
  assign valid_85_io_enable = 1'h0;
  assign valid_85_clock = clock;
  assign valid_85_reset = reset;
  assign valid_86_io_in = 1'h1;
  assign valid_86_io_enable = 1'h0;
  assign valid_86_clock = clock;
  assign valid_86_reset = reset;
  assign valid_87_io_in = 1'h1;
  assign valid_87_io_enable = 1'h0;
  assign valid_87_clock = clock;
  assign valid_87_reset = reset;
  assign valid_88_io_in = 1'h1;
  assign valid_88_io_enable = 1'h0;
  assign valid_88_clock = clock;
  assign valid_88_reset = reset;
  assign valid_89_io_in = 1'h1;
  assign valid_89_io_enable = 1'h0;
  assign valid_89_clock = clock;
  assign valid_89_reset = reset;
  assign valid_90_io_in = 1'h1;
  assign valid_90_io_enable = 1'h0;
  assign valid_90_clock = clock;
  assign valid_90_reset = reset;
  assign valid_91_io_in = 1'h1;
  assign valid_91_io_enable = 1'h0;
  assign valid_91_clock = clock;
  assign valid_91_reset = reset;
  assign valid_92_io_in = 1'h1;
  assign valid_92_io_enable = 1'h0;
  assign valid_92_clock = clock;
  assign valid_92_reset = reset;
  assign valid_93_io_in = 1'h1;
  assign valid_93_io_enable = 1'h0;
  assign valid_93_clock = clock;
  assign valid_93_reset = reset;
  assign valid_94_io_in = 1'h1;
  assign valid_94_io_enable = 1'h0;
  assign valid_94_clock = clock;
  assign valid_94_reset = reset;
  assign valid_95_io_in = 1'h1;
  assign valid_95_io_enable = 1'h0;
  assign valid_95_clock = clock;
  assign valid_95_reset = reset;
  assign valid_96_io_in = 1'h1;
  assign valid_96_io_enable = 1'h0;
  assign valid_96_clock = clock;
  assign valid_96_reset = reset;
  assign valid_97_io_in = 1'h1;
  assign valid_97_io_enable = 1'h0;
  assign valid_97_clock = clock;
  assign valid_97_reset = reset;
  assign valid_98_io_in = 1'h1;
  assign valid_98_io_enable = 1'h0;
  assign valid_98_clock = clock;
  assign valid_98_reset = reset;
  assign valid_99_io_in = 1'h1;
  assign valid_99_io_enable = 1'h0;
  assign valid_99_clock = clock;
  assign valid_99_reset = reset;
  assign valid_100_io_in = 1'h1;
  assign valid_100_io_enable = 1'h0;
  assign valid_100_clock = clock;
  assign valid_100_reset = reset;
  assign valid_101_io_in = 1'h1;
  assign valid_101_io_enable = 1'h0;
  assign valid_101_clock = clock;
  assign valid_101_reset = reset;
  assign valid_102_io_in = 1'h1;
  assign valid_102_io_enable = 1'h0;
  assign valid_102_clock = clock;
  assign valid_102_reset = reset;
  assign valid_103_io_in = 1'h1;
  assign valid_103_io_enable = 1'h0;
  assign valid_103_clock = clock;
  assign valid_103_reset = reset;
  assign valid_104_io_in = 1'h1;
  assign valid_104_io_enable = 1'h0;
  assign valid_104_clock = clock;
  assign valid_104_reset = reset;
  assign valid_105_io_in = 1'h1;
  assign valid_105_io_enable = 1'h0;
  assign valid_105_clock = clock;
  assign valid_105_reset = reset;
  assign valid_106_io_in = 1'h1;
  assign valid_106_io_enable = 1'h0;
  assign valid_106_clock = clock;
  assign valid_106_reset = reset;
  assign valid_107_io_in = 1'h1;
  assign valid_107_io_enable = 1'h0;
  assign valid_107_clock = clock;
  assign valid_107_reset = reset;
  assign valid_108_io_in = 1'h1;
  assign valid_108_io_enable = 1'h0;
  assign valid_108_clock = clock;
  assign valid_108_reset = reset;
  assign valid_109_io_in = 1'h1;
  assign valid_109_io_enable = 1'h0;
  assign valid_109_clock = clock;
  assign valid_109_reset = reset;
  assign valid_110_io_in = 1'h1;
  assign valid_110_io_enable = 1'h0;
  assign valid_110_clock = clock;
  assign valid_110_reset = reset;
  assign valid_111_io_in = 1'h1;
  assign valid_111_io_enable = 1'h0;
  assign valid_111_clock = clock;
  assign valid_111_reset = reset;
  assign valid_112_io_in = 1'h1;
  assign valid_112_io_enable = 1'h0;
  assign valid_112_clock = clock;
  assign valid_112_reset = reset;
  assign valid_113_io_in = 1'h1;
  assign valid_113_io_enable = 1'h0;
  assign valid_113_clock = clock;
  assign valid_113_reset = reset;
  assign valid_114_io_in = 1'h1;
  assign valid_114_io_enable = 1'h0;
  assign valid_114_clock = clock;
  assign valid_114_reset = reset;
  assign valid_115_io_in = 1'h1;
  assign valid_115_io_enable = 1'h0;
  assign valid_115_clock = clock;
  assign valid_115_reset = reset;
  assign valid_116_io_in = 1'h1;
  assign valid_116_io_enable = 1'h0;
  assign valid_116_clock = clock;
  assign valid_116_reset = reset;
  assign valid_117_io_in = 1'h1;
  assign valid_117_io_enable = 1'h0;
  assign valid_117_clock = clock;
  assign valid_117_reset = reset;
  assign valid_118_io_in = 1'h1;
  assign valid_118_io_enable = 1'h0;
  assign valid_118_clock = clock;
  assign valid_118_reset = reset;
  assign valid_119_io_in = 1'h1;
  assign valid_119_io_enable = 1'h0;
  assign valid_119_clock = clock;
  assign valid_119_reset = reset;
  assign valid_120_io_in = 1'h1;
  assign valid_120_io_enable = 1'h0;
  assign valid_120_clock = clock;
  assign valid_120_reset = reset;
  assign valid_121_io_in = 1'h1;
  assign valid_121_io_enable = 1'h0;
  assign valid_121_clock = clock;
  assign valid_121_reset = reset;
  assign valid_122_io_in = 1'h1;
  assign valid_122_io_enable = 1'h0;
  assign valid_122_clock = clock;
  assign valid_122_reset = reset;
  assign valid_123_io_in = 1'h1;
  assign valid_123_io_enable = 1'h0;
  assign valid_123_clock = clock;
  assign valid_123_reset = reset;
  assign valid_124_io_in = 1'h1;
  assign valid_124_io_enable = 1'h0;
  assign valid_124_clock = clock;
  assign valid_124_reset = reset;
  assign valid_125_io_in = 1'h1;
  assign valid_125_io_enable = 1'h0;
  assign valid_125_clock = clock;
  assign valid_125_reset = reset;
  assign valid_126_io_in = 1'h1;
  assign valid_126_io_enable = 1'h0;
  assign valid_126_clock = clock;
  assign valid_126_reset = reset;
  assign valid_127_io_in = 1'h1;
  assign valid_127_io_enable = 1'h0;
  assign valid_127_clock = clock;
  assign valid_127_reset = reset;
  assign valid_128_io_in = 1'h1;
  assign valid_128_io_enable = 1'h0;
  assign valid_128_clock = clock;
  assign valid_128_reset = reset;
  assign valid_129_io_in = 1'h1;
  assign valid_129_io_enable = 1'h0;
  assign valid_129_clock = clock;
  assign valid_129_reset = reset;
  assign valid_130_io_in = 1'h1;
  assign valid_130_io_enable = 1'h0;
  assign valid_130_clock = clock;
  assign valid_130_reset = reset;
  assign valid_131_io_in = 1'h1;
  assign valid_131_io_enable = 1'h0;
  assign valid_131_clock = clock;
  assign valid_131_reset = reset;
  assign valid_132_io_in = 1'h1;
  assign valid_132_io_enable = 1'h0;
  assign valid_132_clock = clock;
  assign valid_132_reset = reset;
  assign valid_133_io_in = 1'h1;
  assign valid_133_io_enable = 1'h0;
  assign valid_133_clock = clock;
  assign valid_133_reset = reset;
  assign valid_134_io_in = 1'h1;
  assign valid_134_io_enable = 1'h0;
  assign valid_134_clock = clock;
  assign valid_134_reset = reset;
  assign valid_135_io_in = 1'h1;
  assign valid_135_io_enable = 1'h0;
  assign valid_135_clock = clock;
  assign valid_135_reset = reset;
  assign valid_136_io_in = 1'h1;
  assign valid_136_io_enable = 1'h0;
  assign valid_136_clock = clock;
  assign valid_136_reset = reset;
  assign valid_137_io_in = 1'h1;
  assign valid_137_io_enable = 1'h0;
  assign valid_137_clock = clock;
  assign valid_137_reset = reset;
  assign valid_138_io_in = 1'h1;
  assign valid_138_io_enable = 1'h0;
  assign valid_138_clock = clock;
  assign valid_138_reset = reset;
  assign valid_139_io_in = 1'h1;
  assign valid_139_io_enable = 1'h0;
  assign valid_139_clock = clock;
  assign valid_139_reset = reset;
  assign valid_140_io_in = 1'h1;
  assign valid_140_io_enable = 1'h0;
  assign valid_140_clock = clock;
  assign valid_140_reset = reset;
  assign valid_141_io_in = 1'h1;
  assign valid_141_io_enable = 1'h0;
  assign valid_141_clock = clock;
  assign valid_141_reset = reset;
  assign valid_142_io_in = 1'h1;
  assign valid_142_io_enable = 1'h0;
  assign valid_142_clock = clock;
  assign valid_142_reset = reset;
  assign valid_143_io_in = 1'h1;
  assign valid_143_io_enable = 1'h0;
  assign valid_143_clock = clock;
  assign valid_143_reset = reset;
  assign valid_144_io_in = 1'h1;
  assign valid_144_io_enable = 1'h0;
  assign valid_144_clock = clock;
  assign valid_144_reset = reset;
  assign valid_145_io_in = 1'h1;
  assign valid_145_io_enable = 1'h0;
  assign valid_145_clock = clock;
  assign valid_145_reset = reset;
  assign valid_146_io_in = 1'h1;
  assign valid_146_io_enable = 1'h0;
  assign valid_146_clock = clock;
  assign valid_146_reset = reset;
  assign valid_147_io_in = 1'h1;
  assign valid_147_io_enable = 1'h0;
  assign valid_147_clock = clock;
  assign valid_147_reset = reset;
  assign valid_148_io_in = 1'h1;
  assign valid_148_io_enable = 1'h0;
  assign valid_148_clock = clock;
  assign valid_148_reset = reset;
  assign valid_149_io_in = 1'h1;
  assign valid_149_io_enable = 1'h0;
  assign valid_149_clock = clock;
  assign valid_149_reset = reset;
  assign valid_150_io_in = 1'h1;
  assign valid_150_io_enable = 1'h0;
  assign valid_150_clock = clock;
  assign valid_150_reset = reset;
  assign valid_151_io_in = 1'h1;
  assign valid_151_io_enable = 1'h0;
  assign valid_151_clock = clock;
  assign valid_151_reset = reset;
  assign valid_152_io_in = 1'h1;
  assign valid_152_io_enable = 1'h0;
  assign valid_152_clock = clock;
  assign valid_152_reset = reset;
  assign valid_153_io_in = 1'h1;
  assign valid_153_io_enable = 1'h0;
  assign valid_153_clock = clock;
  assign valid_153_reset = reset;
  assign valid_154_io_in = 1'h1;
  assign valid_154_io_enable = 1'h0;
  assign valid_154_clock = clock;
  assign valid_154_reset = reset;
  assign valid_155_io_in = 1'h1;
  assign valid_155_io_enable = 1'h0;
  assign valid_155_clock = clock;
  assign valid_155_reset = reset;
  assign valid_156_io_in = 1'h1;
  assign valid_156_io_enable = 1'h0;
  assign valid_156_clock = clock;
  assign valid_156_reset = reset;
  assign valid_157_io_in = 1'h1;
  assign valid_157_io_enable = 1'h0;
  assign valid_157_clock = clock;
  assign valid_157_reset = reset;
  assign valid_158_io_in = 1'h1;
  assign valid_158_io_enable = 1'h0;
  assign valid_158_clock = clock;
  assign valid_158_reset = reset;
  assign valid_159_io_in = 1'h1;
  assign valid_159_io_enable = 1'h0;
  assign valid_159_clock = clock;
  assign valid_159_reset = reset;
  assign valid_160_io_in = 1'h1;
  assign valid_160_io_enable = 1'h0;
  assign valid_160_clock = clock;
  assign valid_160_reset = reset;
  assign valid_161_io_in = 1'h1;
  assign valid_161_io_enable = 1'h0;
  assign valid_161_clock = clock;
  assign valid_161_reset = reset;
  assign valid_162_io_in = 1'h1;
  assign valid_162_io_enable = 1'h0;
  assign valid_162_clock = clock;
  assign valid_162_reset = reset;
  assign valid_163_io_in = 1'h1;
  assign valid_163_io_enable = 1'h0;
  assign valid_163_clock = clock;
  assign valid_163_reset = reset;
  assign valid_164_io_in = 1'h1;
  assign valid_164_io_enable = 1'h0;
  assign valid_164_clock = clock;
  assign valid_164_reset = reset;
  assign valid_165_io_in = 1'h1;
  assign valid_165_io_enable = 1'h0;
  assign valid_165_clock = clock;
  assign valid_165_reset = reset;
  assign valid_166_io_in = 1'h1;
  assign valid_166_io_enable = 1'h0;
  assign valid_166_clock = clock;
  assign valid_166_reset = reset;
  assign valid_167_io_in = 1'h1;
  assign valid_167_io_enable = 1'h0;
  assign valid_167_clock = clock;
  assign valid_167_reset = reset;
  assign valid_168_io_in = 1'h1;
  assign valid_168_io_enable = 1'h0;
  assign valid_168_clock = clock;
  assign valid_168_reset = reset;
  assign valid_169_io_in = 1'h1;
  assign valid_169_io_enable = 1'h0;
  assign valid_169_clock = clock;
  assign valid_169_reset = reset;
  assign valid_170_io_in = 1'h1;
  assign valid_170_io_enable = 1'h0;
  assign valid_170_clock = clock;
  assign valid_170_reset = reset;
  assign valid_171_io_in = 1'h1;
  assign valid_171_io_enable = 1'h0;
  assign valid_171_clock = clock;
  assign valid_171_reset = reset;
  assign valid_172_io_in = 1'h1;
  assign valid_172_io_enable = 1'h0;
  assign valid_172_clock = clock;
  assign valid_172_reset = reset;
  assign valid_173_io_in = 1'h1;
  assign valid_173_io_enable = 1'h0;
  assign valid_173_clock = clock;
  assign valid_173_reset = reset;
  assign valid_174_io_in = 1'h1;
  assign valid_174_io_enable = 1'h0;
  assign valid_174_clock = clock;
  assign valid_174_reset = reset;
  assign valid_175_io_in = 1'h1;
  assign valid_175_io_enable = 1'h0;
  assign valid_175_clock = clock;
  assign valid_175_reset = reset;
  assign valid_176_io_in = 1'h1;
  assign valid_176_io_enable = 1'h0;
  assign valid_176_clock = clock;
  assign valid_176_reset = reset;
  assign valid_177_io_in = 1'h1;
  assign valid_177_io_enable = 1'h0;
  assign valid_177_clock = clock;
  assign valid_177_reset = reset;
  assign valid_178_io_in = 1'h1;
  assign valid_178_io_enable = 1'h0;
  assign valid_178_clock = clock;
  assign valid_178_reset = reset;
  assign valid_179_io_in = 1'h1;
  assign valid_179_io_enable = 1'h0;
  assign valid_179_clock = clock;
  assign valid_179_reset = reset;
  assign valid_180_io_in = 1'h1;
  assign valid_180_io_enable = 1'h0;
  assign valid_180_clock = clock;
  assign valid_180_reset = reset;
  assign valid_181_io_in = 1'h1;
  assign valid_181_io_enable = 1'h0;
  assign valid_181_clock = clock;
  assign valid_181_reset = reset;
  assign valid_182_io_in = 1'h1;
  assign valid_182_io_enable = 1'h0;
  assign valid_182_clock = clock;
  assign valid_182_reset = reset;
  assign valid_183_io_in = 1'h1;
  assign valid_183_io_enable = 1'h0;
  assign valid_183_clock = clock;
  assign valid_183_reset = reset;
  assign valid_184_io_in = 1'h1;
  assign valid_184_io_enable = 1'h0;
  assign valid_184_clock = clock;
  assign valid_184_reset = reset;
  assign valid_185_io_in = 1'h1;
  assign valid_185_io_enable = 1'h0;
  assign valid_185_clock = clock;
  assign valid_185_reset = reset;
  assign valid_186_io_in = 1'h1;
  assign valid_186_io_enable = 1'h0;
  assign valid_186_clock = clock;
  assign valid_186_reset = reset;
  assign valid_187_io_in = 1'h1;
  assign valid_187_io_enable = 1'h0;
  assign valid_187_clock = clock;
  assign valid_187_reset = reset;
  assign valid_188_io_in = 1'h1;
  assign valid_188_io_enable = 1'h0;
  assign valid_188_clock = clock;
  assign valid_188_reset = reset;
  assign valid_189_io_in = 1'h1;
  assign valid_189_io_enable = 1'h0;
  assign valid_189_clock = clock;
  assign valid_189_reset = reset;
  assign valid_190_io_in = 1'h1;
  assign valid_190_io_enable = 1'h0;
  assign valid_190_clock = clock;
  assign valid_190_reset = reset;
  assign valid_191_io_in = 1'h1;
  assign valid_191_io_enable = 1'h0;
  assign valid_191_clock = clock;
  assign valid_191_reset = reset;
  assign valid_192_io_in = 1'h1;
  assign valid_192_io_enable = 1'h0;
  assign valid_192_clock = clock;
  assign valid_192_reset = reset;
  assign valid_193_io_in = 1'h1;
  assign valid_193_io_enable = 1'h0;
  assign valid_193_clock = clock;
  assign valid_193_reset = reset;
  assign valid_194_io_in = 1'h1;
  assign valid_194_io_enable = 1'h0;
  assign valid_194_clock = clock;
  assign valid_194_reset = reset;
  assign valid_195_io_in = 1'h1;
  assign valid_195_io_enable = 1'h0;
  assign valid_195_clock = clock;
  assign valid_195_reset = reset;
  assign valid_196_io_in = 1'h1;
  assign valid_196_io_enable = 1'h0;
  assign valid_196_clock = clock;
  assign valid_196_reset = reset;
  assign valid_197_io_in = 1'h1;
  assign valid_197_io_enable = 1'h0;
  assign valid_197_clock = clock;
  assign valid_197_reset = reset;
  assign valid_198_io_in = 1'h1;
  assign valid_198_io_enable = 1'h0;
  assign valid_198_clock = clock;
  assign valid_198_reset = reset;
  assign valid_199_io_in = 1'h1;
  assign valid_199_io_enable = 1'h0;
  assign valid_199_clock = clock;
  assign valid_199_reset = reset;
  assign valid_200_io_in = 1'h1;
  assign valid_200_io_enable = 1'h0;
  assign valid_200_clock = clock;
  assign valid_200_reset = reset;
  assign valid_201_io_in = 1'h1;
  assign valid_201_io_enable = 1'h0;
  assign valid_201_clock = clock;
  assign valid_201_reset = reset;
  assign valid_202_io_in = 1'h1;
  assign valid_202_io_enable = 1'h0;
  assign valid_202_clock = clock;
  assign valid_202_reset = reset;
  assign valid_203_io_in = 1'h1;
  assign valid_203_io_enable = 1'h0;
  assign valid_203_clock = clock;
  assign valid_203_reset = reset;
  assign valid_204_io_in = 1'h1;
  assign valid_204_io_enable = 1'h0;
  assign valid_204_clock = clock;
  assign valid_204_reset = reset;
  assign valid_205_io_in = 1'h1;
  assign valid_205_io_enable = 1'h0;
  assign valid_205_clock = clock;
  assign valid_205_reset = reset;
  assign valid_206_io_in = 1'h1;
  assign valid_206_io_enable = 1'h0;
  assign valid_206_clock = clock;
  assign valid_206_reset = reset;
  assign valid_207_io_in = 1'h1;
  assign valid_207_io_enable = 1'h0;
  assign valid_207_clock = clock;
  assign valid_207_reset = reset;
  assign valid_208_io_in = 1'h1;
  assign valid_208_io_enable = 1'h0;
  assign valid_208_clock = clock;
  assign valid_208_reset = reset;
  assign valid_209_io_in = 1'h1;
  assign valid_209_io_enable = 1'h0;
  assign valid_209_clock = clock;
  assign valid_209_reset = reset;
  assign valid_210_io_in = 1'h1;
  assign valid_210_io_enable = 1'h0;
  assign valid_210_clock = clock;
  assign valid_210_reset = reset;
  assign valid_211_io_in = 1'h1;
  assign valid_211_io_enable = 1'h0;
  assign valid_211_clock = clock;
  assign valid_211_reset = reset;
  assign valid_212_io_in = 1'h1;
  assign valid_212_io_enable = 1'h0;
  assign valid_212_clock = clock;
  assign valid_212_reset = reset;
  assign valid_213_io_in = 1'h1;
  assign valid_213_io_enable = 1'h0;
  assign valid_213_clock = clock;
  assign valid_213_reset = reset;
  assign valid_214_io_in = 1'h1;
  assign valid_214_io_enable = 1'h0;
  assign valid_214_clock = clock;
  assign valid_214_reset = reset;
  assign valid_215_io_in = 1'h1;
  assign valid_215_io_enable = 1'h0;
  assign valid_215_clock = clock;
  assign valid_215_reset = reset;
  assign valid_216_io_in = 1'h1;
  assign valid_216_io_enable = 1'h0;
  assign valid_216_clock = clock;
  assign valid_216_reset = reset;
  assign valid_217_io_in = 1'h1;
  assign valid_217_io_enable = 1'h0;
  assign valid_217_clock = clock;
  assign valid_217_reset = reset;
  assign valid_218_io_in = 1'h1;
  assign valid_218_io_enable = 1'h0;
  assign valid_218_clock = clock;
  assign valid_218_reset = reset;
  assign valid_219_io_in = 1'h1;
  assign valid_219_io_enable = 1'h0;
  assign valid_219_clock = clock;
  assign valid_219_reset = reset;
  assign valid_220_io_in = 1'h1;
  assign valid_220_io_enable = 1'h0;
  assign valid_220_clock = clock;
  assign valid_220_reset = reset;
  assign valid_221_io_in = 1'h1;
  assign valid_221_io_enable = 1'h0;
  assign valid_221_clock = clock;
  assign valid_221_reset = reset;
  assign valid_222_io_in = 1'h1;
  assign valid_222_io_enable = 1'h0;
  assign valid_222_clock = clock;
  assign valid_222_reset = reset;
  assign valid_223_io_in = 1'h1;
  assign valid_223_io_enable = 1'h0;
  assign valid_223_clock = clock;
  assign valid_223_reset = reset;
  assign valid_224_io_in = 1'h1;
  assign valid_224_io_enable = 1'h0;
  assign valid_224_clock = clock;
  assign valid_224_reset = reset;
  assign valid_225_io_in = 1'h1;
  assign valid_225_io_enable = 1'h0;
  assign valid_225_clock = clock;
  assign valid_225_reset = reset;
  assign valid_226_io_in = 1'h1;
  assign valid_226_io_enable = 1'h0;
  assign valid_226_clock = clock;
  assign valid_226_reset = reset;
  assign valid_227_io_in = 1'h1;
  assign valid_227_io_enable = 1'h0;
  assign valid_227_clock = clock;
  assign valid_227_reset = reset;
  assign valid_228_io_in = 1'h1;
  assign valid_228_io_enable = 1'h0;
  assign valid_228_clock = clock;
  assign valid_228_reset = reset;
  assign valid_229_io_in = 1'h1;
  assign valid_229_io_enable = 1'h0;
  assign valid_229_clock = clock;
  assign valid_229_reset = reset;
  assign valid_230_io_in = 1'h1;
  assign valid_230_io_enable = 1'h0;
  assign valid_230_clock = clock;
  assign valid_230_reset = reset;
  assign valid_231_io_in = 1'h1;
  assign valid_231_io_enable = 1'h0;
  assign valid_231_clock = clock;
  assign valid_231_reset = reset;
  assign valid_232_io_in = 1'h1;
  assign valid_232_io_enable = 1'h0;
  assign valid_232_clock = clock;
  assign valid_232_reset = reset;
  assign valid_233_io_in = 1'h1;
  assign valid_233_io_enable = 1'h0;
  assign valid_233_clock = clock;
  assign valid_233_reset = reset;
  assign valid_234_io_in = 1'h1;
  assign valid_234_io_enable = 1'h0;
  assign valid_234_clock = clock;
  assign valid_234_reset = reset;
  assign valid_235_io_in = 1'h1;
  assign valid_235_io_enable = 1'h0;
  assign valid_235_clock = clock;
  assign valid_235_reset = reset;
  assign valid_236_io_in = 1'h1;
  assign valid_236_io_enable = 1'h0;
  assign valid_236_clock = clock;
  assign valid_236_reset = reset;
  assign valid_237_io_in = 1'h1;
  assign valid_237_io_enable = 1'h0;
  assign valid_237_clock = clock;
  assign valid_237_reset = reset;
  assign valid_238_io_in = 1'h1;
  assign valid_238_io_enable = 1'h0;
  assign valid_238_clock = clock;
  assign valid_238_reset = reset;
  assign valid_239_io_in = 1'h1;
  assign valid_239_io_enable = 1'h0;
  assign valid_239_clock = clock;
  assign valid_239_reset = reset;
  assign valid_240_io_in = 1'h1;
  assign valid_240_io_enable = 1'h0;
  assign valid_240_clock = clock;
  assign valid_240_reset = reset;
  assign valid_241_io_in = 1'h1;
  assign valid_241_io_enable = 1'h0;
  assign valid_241_clock = clock;
  assign valid_241_reset = reset;
  assign valid_242_io_in = 1'h1;
  assign valid_242_io_enable = 1'h0;
  assign valid_242_clock = clock;
  assign valid_242_reset = reset;
  assign valid_243_io_in = 1'h1;
  assign valid_243_io_enable = 1'h0;
  assign valid_243_clock = clock;
  assign valid_243_reset = reset;
  assign valid_244_io_in = 1'h1;
  assign valid_244_io_enable = 1'h0;
  assign valid_244_clock = clock;
  assign valid_244_reset = reset;
  assign valid_245_io_in = 1'h1;
  assign valid_245_io_enable = 1'h0;
  assign valid_245_clock = clock;
  assign valid_245_reset = reset;
  assign valid_246_io_in = 1'h1;
  assign valid_246_io_enable = 1'h0;
  assign valid_246_clock = clock;
  assign valid_246_reset = reset;
  assign valid_247_io_in = 1'h1;
  assign valid_247_io_enable = 1'h0;
  assign valid_247_clock = clock;
  assign valid_247_reset = reset;
  assign valid_248_io_in = 1'h1;
  assign valid_248_io_enable = 1'h0;
  assign valid_248_clock = clock;
  assign valid_248_reset = reset;
  assign valid_249_io_in = 1'h1;
  assign valid_249_io_enable = 1'h0;
  assign valid_249_clock = clock;
  assign valid_249_reset = reset;
  assign valid_250_io_in = 1'h1;
  assign valid_250_io_enable = 1'h0;
  assign valid_250_clock = clock;
  assign valid_250_reset = reset;
  assign valid_251_io_in = 1'h1;
  assign valid_251_io_enable = 1'h0;
  assign valid_251_clock = clock;
  assign valid_251_reset = reset;
  assign valid_252_io_in = 1'h1;
  assign valid_252_io_enable = 1'h0;
  assign valid_252_clock = clock;
  assign valid_252_reset = reset;
  assign valid_253_io_in = 1'h1;
  assign valid_253_io_enable = 1'h0;
  assign valid_253_clock = clock;
  assign valid_253_reset = reset;
  assign valid_254_io_in = 1'h1;
  assign valid_254_io_enable = 1'h0;
  assign valid_254_clock = clock;
  assign valid_254_reset = reset;
  assign valid_255_io_in = 1'h1;
  assign valid_255_io_enable = 1'h0;
  assign valid_255_clock = clock;
  assign valid_255_reset = reset;
  assign valid_256_io_in = 1'h1;
  assign valid_256_io_enable = 1'h0;
  assign valid_256_clock = clock;
  assign valid_256_reset = reset;
  assign valid_257_io_in = 1'h1;
  assign valid_257_io_enable = 1'h0;
  assign valid_257_clock = clock;
  assign valid_257_reset = reset;
  assign valid_258_io_in = 1'h1;
  assign valid_258_io_enable = 1'h0;
  assign valid_258_clock = clock;
  assign valid_258_reset = reset;
  assign valid_259_io_in = 1'h1;
  assign valid_259_io_enable = 1'h0;
  assign valid_259_clock = clock;
  assign valid_259_reset = reset;
  assign valid_260_io_in = 1'h1;
  assign valid_260_io_enable = 1'h0;
  assign valid_260_clock = clock;
  assign valid_260_reset = reset;
  assign valid_261_io_in = 1'h1;
  assign valid_261_io_enable = 1'h0;
  assign valid_261_clock = clock;
  assign valid_261_reset = reset;
  assign valid_262_io_in = 1'h1;
  assign valid_262_io_enable = 1'h0;
  assign valid_262_clock = clock;
  assign valid_262_reset = reset;
  assign valid_263_io_in = 1'h1;
  assign valid_263_io_enable = 1'h0;
  assign valid_263_clock = clock;
  assign valid_263_reset = reset;
  assign valid_264_io_in = 1'h1;
  assign valid_264_io_enable = 1'h0;
  assign valid_264_clock = clock;
  assign valid_264_reset = reset;
  assign valid_265_io_in = 1'h1;
  assign valid_265_io_enable = 1'h0;
  assign valid_265_clock = clock;
  assign valid_265_reset = reset;
  assign valid_266_io_in = 1'h1;
  assign valid_266_io_enable = 1'h0;
  assign valid_266_clock = clock;
  assign valid_266_reset = reset;
  assign valid_267_io_in = 1'h1;
  assign valid_267_io_enable = 1'h0;
  assign valid_267_clock = clock;
  assign valid_267_reset = reset;
  assign valid_268_io_in = 1'h1;
  assign valid_268_io_enable = 1'h0;
  assign valid_268_clock = clock;
  assign valid_268_reset = reset;
  assign valid_269_io_in = 1'h1;
  assign valid_269_io_enable = 1'h0;
  assign valid_269_clock = clock;
  assign valid_269_reset = reset;
  assign valid_270_io_in = 1'h1;
  assign valid_270_io_enable = 1'h0;
  assign valid_270_clock = clock;
  assign valid_270_reset = reset;
  assign valid_271_io_in = 1'h1;
  assign valid_271_io_enable = 1'h0;
  assign valid_271_clock = clock;
  assign valid_271_reset = reset;
  assign valid_272_io_in = 1'h1;
  assign valid_272_io_enable = 1'h0;
  assign valid_272_clock = clock;
  assign valid_272_reset = reset;
  assign valid_273_io_in = 1'h1;
  assign valid_273_io_enable = 1'h0;
  assign valid_273_clock = clock;
  assign valid_273_reset = reset;
  assign valid_274_io_in = 1'h1;
  assign valid_274_io_enable = 1'h0;
  assign valid_274_clock = clock;
  assign valid_274_reset = reset;
  assign valid_275_io_in = 1'h1;
  assign valid_275_io_enable = 1'h0;
  assign valid_275_clock = clock;
  assign valid_275_reset = reset;
  assign valid_276_io_in = 1'h1;
  assign valid_276_io_enable = 1'h0;
  assign valid_276_clock = clock;
  assign valid_276_reset = reset;
  assign valid_277_io_in = 1'h1;
  assign valid_277_io_enable = 1'h0;
  assign valid_277_clock = clock;
  assign valid_277_reset = reset;
  assign valid_278_io_in = 1'h1;
  assign valid_278_io_enable = 1'h0;
  assign valid_278_clock = clock;
  assign valid_278_reset = reset;
  assign valid_279_io_in = 1'h1;
  assign valid_279_io_enable = 1'h0;
  assign valid_279_clock = clock;
  assign valid_279_reset = reset;
  assign valid_280_io_in = 1'h1;
  assign valid_280_io_enable = 1'h0;
  assign valid_280_clock = clock;
  assign valid_280_reset = reset;
  assign valid_281_io_in = 1'h1;
  assign valid_281_io_enable = 1'h0;
  assign valid_281_clock = clock;
  assign valid_281_reset = reset;
  assign valid_282_io_in = 1'h1;
  assign valid_282_io_enable = 1'h0;
  assign valid_282_clock = clock;
  assign valid_282_reset = reset;
  assign valid_283_io_in = 1'h1;
  assign valid_283_io_enable = 1'h0;
  assign valid_283_clock = clock;
  assign valid_283_reset = reset;
  assign valid_284_io_in = 1'h1;
  assign valid_284_io_enable = 1'h0;
  assign valid_284_clock = clock;
  assign valid_284_reset = reset;
  assign valid_285_io_in = 1'h1;
  assign valid_285_io_enable = 1'h0;
  assign valid_285_clock = clock;
  assign valid_285_reset = reset;
  assign valid_286_io_in = 1'h1;
  assign valid_286_io_enable = 1'h0;
  assign valid_286_clock = clock;
  assign valid_286_reset = reset;
  assign valid_287_io_in = 1'h1;
  assign valid_287_io_enable = 1'h0;
  assign valid_287_clock = clock;
  assign valid_287_reset = reset;
  assign valid_288_io_in = 1'h1;
  assign valid_288_io_enable = 1'h0;
  assign valid_288_clock = clock;
  assign valid_288_reset = reset;
  assign valid_289_io_in = 1'h1;
  assign valid_289_io_enable = 1'h0;
  assign valid_289_clock = clock;
  assign valid_289_reset = reset;
  assign valid_290_io_in = 1'h1;
  assign valid_290_io_enable = 1'h0;
  assign valid_290_clock = clock;
  assign valid_290_reset = reset;
  assign valid_291_io_in = 1'h1;
  assign valid_291_io_enable = 1'h0;
  assign valid_291_clock = clock;
  assign valid_291_reset = reset;
  assign valid_292_io_in = 1'h1;
  assign valid_292_io_enable = 1'h0;
  assign valid_292_clock = clock;
  assign valid_292_reset = reset;
  assign valid_293_io_in = 1'h1;
  assign valid_293_io_enable = 1'h0;
  assign valid_293_clock = clock;
  assign valid_293_reset = reset;
  assign valid_294_io_in = 1'h1;
  assign valid_294_io_enable = 1'h0;
  assign valid_294_clock = clock;
  assign valid_294_reset = reset;
  assign valid_295_io_in = 1'h1;
  assign valid_295_io_enable = 1'h0;
  assign valid_295_clock = clock;
  assign valid_295_reset = reset;
  assign valid_296_io_in = 1'h1;
  assign valid_296_io_enable = 1'h0;
  assign valid_296_clock = clock;
  assign valid_296_reset = reset;
  assign valid_297_io_in = 1'h1;
  assign valid_297_io_enable = 1'h0;
  assign valid_297_clock = clock;
  assign valid_297_reset = reset;
  assign valid_298_io_in = 1'h1;
  assign valid_298_io_enable = 1'h0;
  assign valid_298_clock = clock;
  assign valid_298_reset = reset;
  assign valid_299_io_in = 1'h1;
  assign valid_299_io_enable = 1'h0;
  assign valid_299_clock = clock;
  assign valid_299_reset = reset;
  assign valid_300_io_in = 1'h1;
  assign valid_300_io_enable = 1'h0;
  assign valid_300_clock = clock;
  assign valid_300_reset = reset;
  assign valid_301_io_in = 1'h1;
  assign valid_301_io_enable = 1'h0;
  assign valid_301_clock = clock;
  assign valid_301_reset = reset;
  assign valid_302_io_in = 1'h1;
  assign valid_302_io_enable = 1'h0;
  assign valid_302_clock = clock;
  assign valid_302_reset = reset;
  assign valid_303_io_in = 1'h1;
  assign valid_303_io_enable = 1'h0;
  assign valid_303_clock = clock;
  assign valid_303_reset = reset;
  assign valid_304_io_in = 1'h1;
  assign valid_304_io_enable = 1'h0;
  assign valid_304_clock = clock;
  assign valid_304_reset = reset;
  assign valid_305_io_in = 1'h1;
  assign valid_305_io_enable = 1'h0;
  assign valid_305_clock = clock;
  assign valid_305_reset = reset;
  assign valid_306_io_in = 1'h1;
  assign valid_306_io_enable = 1'h0;
  assign valid_306_clock = clock;
  assign valid_306_reset = reset;
  assign valid_307_io_in = 1'h1;
  assign valid_307_io_enable = 1'h0;
  assign valid_307_clock = clock;
  assign valid_307_reset = reset;
  assign valid_308_io_in = 1'h1;
  assign valid_308_io_enable = 1'h0;
  assign valid_308_clock = clock;
  assign valid_308_reset = reset;
  assign valid_309_io_in = 1'h1;
  assign valid_309_io_enable = 1'h0;
  assign valid_309_clock = clock;
  assign valid_309_reset = reset;
  assign valid_310_io_in = 1'h1;
  assign valid_310_io_enable = 1'h0;
  assign valid_310_clock = clock;
  assign valid_310_reset = reset;
  assign valid_311_io_in = 1'h1;
  assign valid_311_io_enable = 1'h0;
  assign valid_311_clock = clock;
  assign valid_311_reset = reset;
  assign valid_312_io_in = 1'h1;
  assign valid_312_io_enable = 1'h0;
  assign valid_312_clock = clock;
  assign valid_312_reset = reset;
  assign valid_313_io_in = 1'h1;
  assign valid_313_io_enable = 1'h0;
  assign valid_313_clock = clock;
  assign valid_313_reset = reset;
  assign valid_314_io_in = 1'h1;
  assign valid_314_io_enable = 1'h0;
  assign valid_314_clock = clock;
  assign valid_314_reset = reset;
  assign valid_315_io_in = 1'h1;
  assign valid_315_io_enable = 1'h0;
  assign valid_315_clock = clock;
  assign valid_315_reset = reset;
  assign valid_316_io_in = 1'h1;
  assign valid_316_io_enable = 1'h0;
  assign valid_316_clock = clock;
  assign valid_316_reset = reset;
  assign valid_317_io_in = 1'h1;
  assign valid_317_io_enable = 1'h0;
  assign valid_317_clock = clock;
  assign valid_317_reset = reset;
  assign valid_318_io_in = 1'h1;
  assign valid_318_io_enable = 1'h0;
  assign valid_318_clock = clock;
  assign valid_318_reset = reset;
  assign valid_319_io_in = 1'h1;
  assign valid_319_io_enable = 1'h0;
  assign valid_319_clock = clock;
  assign valid_319_reset = reset;
  assign valid_320_io_in = 1'h1;
  assign valid_320_io_enable = 1'h0;
  assign valid_320_clock = clock;
  assign valid_320_reset = reset;
  assign valid_321_io_in = 1'h1;
  assign valid_321_io_enable = 1'h0;
  assign valid_321_clock = clock;
  assign valid_321_reset = reset;
  assign valid_322_io_in = 1'h1;
  assign valid_322_io_enable = 1'h0;
  assign valid_322_clock = clock;
  assign valid_322_reset = reset;
  assign valid_323_io_in = 1'h1;
  assign valid_323_io_enable = 1'h0;
  assign valid_323_clock = clock;
  assign valid_323_reset = reset;
  assign valid_324_io_in = 1'h1;
  assign valid_324_io_enable = 1'h0;
  assign valid_324_clock = clock;
  assign valid_324_reset = reset;
  assign valid_325_io_in = 1'h1;
  assign valid_325_io_enable = 1'h0;
  assign valid_325_clock = clock;
  assign valid_325_reset = reset;
  assign valid_326_io_in = 1'h1;
  assign valid_326_io_enable = 1'h0;
  assign valid_326_clock = clock;
  assign valid_326_reset = reset;
  assign valid_327_io_in = 1'h1;
  assign valid_327_io_enable = 1'h0;
  assign valid_327_clock = clock;
  assign valid_327_reset = reset;
  assign valid_328_io_in = 1'h1;
  assign valid_328_io_enable = 1'h0;
  assign valid_328_clock = clock;
  assign valid_328_reset = reset;
  assign valid_329_io_in = 1'h1;
  assign valid_329_io_enable = 1'h0;
  assign valid_329_clock = clock;
  assign valid_329_reset = reset;
  assign valid_330_io_in = 1'h1;
  assign valid_330_io_enable = 1'h0;
  assign valid_330_clock = clock;
  assign valid_330_reset = reset;
  assign valid_331_io_in = 1'h1;
  assign valid_331_io_enable = 1'h0;
  assign valid_331_clock = clock;
  assign valid_331_reset = reset;
  assign valid_332_io_in = 1'h1;
  assign valid_332_io_enable = 1'h0;
  assign valid_332_clock = clock;
  assign valid_332_reset = reset;
  assign valid_333_io_in = 1'h1;
  assign valid_333_io_enable = 1'h0;
  assign valid_333_clock = clock;
  assign valid_333_reset = reset;
  assign valid_334_io_in = 1'h1;
  assign valid_334_io_enable = 1'h0;
  assign valid_334_clock = clock;
  assign valid_334_reset = reset;
  assign valid_335_io_in = 1'h1;
  assign valid_335_io_enable = 1'h0;
  assign valid_335_clock = clock;
  assign valid_335_reset = reset;
  assign valid_336_io_in = 1'h1;
  assign valid_336_io_enable = 1'h0;
  assign valid_336_clock = clock;
  assign valid_336_reset = reset;
  assign valid_337_io_in = 1'h1;
  assign valid_337_io_enable = 1'h0;
  assign valid_337_clock = clock;
  assign valid_337_reset = reset;
  assign valid_338_io_in = 1'h1;
  assign valid_338_io_enable = 1'h0;
  assign valid_338_clock = clock;
  assign valid_338_reset = reset;
  assign valid_339_io_in = 1'h1;
  assign valid_339_io_enable = 1'h0;
  assign valid_339_clock = clock;
  assign valid_339_reset = reset;
  assign valid_340_io_in = 1'h1;
  assign valid_340_io_enable = 1'h0;
  assign valid_340_clock = clock;
  assign valid_340_reset = reset;
  assign valid_341_io_in = 1'h1;
  assign valid_341_io_enable = 1'h0;
  assign valid_341_clock = clock;
  assign valid_341_reset = reset;
  assign valid_342_io_in = 1'h1;
  assign valid_342_io_enable = 1'h0;
  assign valid_342_clock = clock;
  assign valid_342_reset = reset;
  assign valid_343_io_in = 1'h1;
  assign valid_343_io_enable = 1'h0;
  assign valid_343_clock = clock;
  assign valid_343_reset = reset;
  assign valid_344_io_in = 1'h1;
  assign valid_344_io_enable = 1'h0;
  assign valid_344_clock = clock;
  assign valid_344_reset = reset;
  assign valid_345_io_in = 1'h1;
  assign valid_345_io_enable = 1'h0;
  assign valid_345_clock = clock;
  assign valid_345_reset = reset;
  assign valid_346_io_in = 1'h1;
  assign valid_346_io_enable = 1'h0;
  assign valid_346_clock = clock;
  assign valid_346_reset = reset;
  assign valid_347_io_in = 1'h1;
  assign valid_347_io_enable = 1'h0;
  assign valid_347_clock = clock;
  assign valid_347_reset = reset;
  assign valid_348_io_in = 1'h1;
  assign valid_348_io_enable = 1'h0;
  assign valid_348_clock = clock;
  assign valid_348_reset = reset;
  assign valid_349_io_in = 1'h1;
  assign valid_349_io_enable = 1'h0;
  assign valid_349_clock = clock;
  assign valid_349_reset = reset;
  assign valid_350_io_in = 1'h1;
  assign valid_350_io_enable = 1'h0;
  assign valid_350_clock = clock;
  assign valid_350_reset = reset;
  assign valid_351_io_in = 1'h1;
  assign valid_351_io_enable = 1'h0;
  assign valid_351_clock = clock;
  assign valid_351_reset = reset;
  assign valid_352_io_in = 1'h1;
  assign valid_352_io_enable = 1'h0;
  assign valid_352_clock = clock;
  assign valid_352_reset = reset;
  assign valid_353_io_in = 1'h1;
  assign valid_353_io_enable = 1'h0;
  assign valid_353_clock = clock;
  assign valid_353_reset = reset;
  assign valid_354_io_in = 1'h1;
  assign valid_354_io_enable = 1'h0;
  assign valid_354_clock = clock;
  assign valid_354_reset = reset;
  assign valid_355_io_in = 1'h1;
  assign valid_355_io_enable = 1'h0;
  assign valid_355_clock = clock;
  assign valid_355_reset = reset;
  assign valid_356_io_in = 1'h1;
  assign valid_356_io_enable = 1'h0;
  assign valid_356_clock = clock;
  assign valid_356_reset = reset;
  assign valid_357_io_in = 1'h1;
  assign valid_357_io_enable = 1'h0;
  assign valid_357_clock = clock;
  assign valid_357_reset = reset;
  assign valid_358_io_in = 1'h1;
  assign valid_358_io_enable = 1'h0;
  assign valid_358_clock = clock;
  assign valid_358_reset = reset;
  assign valid_359_io_in = 1'h1;
  assign valid_359_io_enable = 1'h0;
  assign valid_359_clock = clock;
  assign valid_359_reset = reset;
  assign valid_360_io_in = 1'h1;
  assign valid_360_io_enable = 1'h0;
  assign valid_360_clock = clock;
  assign valid_360_reset = reset;
  assign valid_361_io_in = 1'h1;
  assign valid_361_io_enable = 1'h0;
  assign valid_361_clock = clock;
  assign valid_361_reset = reset;
  assign valid_362_io_in = 1'h1;
  assign valid_362_io_enable = 1'h0;
  assign valid_362_clock = clock;
  assign valid_362_reset = reset;
  assign valid_363_io_in = 1'h1;
  assign valid_363_io_enable = 1'h0;
  assign valid_363_clock = clock;
  assign valid_363_reset = reset;
  assign valid_364_io_in = 1'h1;
  assign valid_364_io_enable = 1'h0;
  assign valid_364_clock = clock;
  assign valid_364_reset = reset;
  assign valid_365_io_in = 1'h1;
  assign valid_365_io_enable = 1'h0;
  assign valid_365_clock = clock;
  assign valid_365_reset = reset;
  assign valid_366_io_in = 1'h1;
  assign valid_366_io_enable = 1'h0;
  assign valid_366_clock = clock;
  assign valid_366_reset = reset;
  assign valid_367_io_in = 1'h1;
  assign valid_367_io_enable = 1'h0;
  assign valid_367_clock = clock;
  assign valid_367_reset = reset;
  assign valid_368_io_in = 1'h1;
  assign valid_368_io_enable = 1'h0;
  assign valid_368_clock = clock;
  assign valid_368_reset = reset;
  assign valid_369_io_in = 1'h1;
  assign valid_369_io_enable = 1'h0;
  assign valid_369_clock = clock;
  assign valid_369_reset = reset;
  assign valid_370_io_in = 1'h1;
  assign valid_370_io_enable = 1'h0;
  assign valid_370_clock = clock;
  assign valid_370_reset = reset;
  assign valid_371_io_in = 1'h1;
  assign valid_371_io_enable = 1'h0;
  assign valid_371_clock = clock;
  assign valid_371_reset = reset;
  assign valid_372_io_in = 1'h1;
  assign valid_372_io_enable = 1'h0;
  assign valid_372_clock = clock;
  assign valid_372_reset = reset;
  assign valid_373_io_in = 1'h1;
  assign valid_373_io_enable = 1'h0;
  assign valid_373_clock = clock;
  assign valid_373_reset = reset;
  assign valid_374_io_in = 1'h1;
  assign valid_374_io_enable = 1'h0;
  assign valid_374_clock = clock;
  assign valid_374_reset = reset;
  assign valid_375_io_in = 1'h1;
  assign valid_375_io_enable = 1'h0;
  assign valid_375_clock = clock;
  assign valid_375_reset = reset;
  assign valid_376_io_in = 1'h1;
  assign valid_376_io_enable = 1'h0;
  assign valid_376_clock = clock;
  assign valid_376_reset = reset;
  assign valid_377_io_in = 1'h1;
  assign valid_377_io_enable = 1'h0;
  assign valid_377_clock = clock;
  assign valid_377_reset = reset;
  assign valid_378_io_in = 1'h1;
  assign valid_378_io_enable = 1'h0;
  assign valid_378_clock = clock;
  assign valid_378_reset = reset;
  assign valid_379_io_in = 1'h1;
  assign valid_379_io_enable = 1'h0;
  assign valid_379_clock = clock;
  assign valid_379_reset = reset;
  assign valid_380_io_in = 1'h1;
  assign valid_380_io_enable = 1'h0;
  assign valid_380_clock = clock;
  assign valid_380_reset = reset;
  assign valid_381_io_in = 1'h1;
  assign valid_381_io_enable = 1'h0;
  assign valid_381_clock = clock;
  assign valid_381_reset = reset;
  assign valid_382_io_in = 1'h1;
  assign valid_382_io_enable = 1'h0;
  assign valid_382_clock = clock;
  assign valid_382_reset = reset;
  assign valid_383_io_in = 1'h1;
  assign valid_383_io_enable = 1'h0;
  assign valid_383_clock = clock;
  assign valid_383_reset = reset;
  assign valid_384_io_in = 1'h1;
  assign valid_384_io_enable = 1'h0;
  assign valid_384_clock = clock;
  assign valid_384_reset = reset;
  assign valid_385_io_in = 1'h1;
  assign valid_385_io_enable = 1'h0;
  assign valid_385_clock = clock;
  assign valid_385_reset = reset;
  assign valid_386_io_in = 1'h1;
  assign valid_386_io_enable = 1'h0;
  assign valid_386_clock = clock;
  assign valid_386_reset = reset;
  assign valid_387_io_in = 1'h1;
  assign valid_387_io_enable = 1'h0;
  assign valid_387_clock = clock;
  assign valid_387_reset = reset;
  assign valid_388_io_in = 1'h1;
  assign valid_388_io_enable = 1'h0;
  assign valid_388_clock = clock;
  assign valid_388_reset = reset;
  assign valid_389_io_in = 1'h1;
  assign valid_389_io_enable = 1'h0;
  assign valid_389_clock = clock;
  assign valid_389_reset = reset;
  assign valid_390_io_in = 1'h1;
  assign valid_390_io_enable = 1'h0;
  assign valid_390_clock = clock;
  assign valid_390_reset = reset;
  assign valid_391_io_in = 1'h1;
  assign valid_391_io_enable = 1'h0;
  assign valid_391_clock = clock;
  assign valid_391_reset = reset;
  assign valid_392_io_in = 1'h1;
  assign valid_392_io_enable = 1'h0;
  assign valid_392_clock = clock;
  assign valid_392_reset = reset;
  assign valid_393_io_in = 1'h1;
  assign valid_393_io_enable = 1'h0;
  assign valid_393_clock = clock;
  assign valid_393_reset = reset;
  assign valid_394_io_in = 1'h1;
  assign valid_394_io_enable = 1'h0;
  assign valid_394_clock = clock;
  assign valid_394_reset = reset;
  assign valid_395_io_in = 1'h1;
  assign valid_395_io_enable = 1'h0;
  assign valid_395_clock = clock;
  assign valid_395_reset = reset;
  assign valid_396_io_in = 1'h1;
  assign valid_396_io_enable = 1'h0;
  assign valid_396_clock = clock;
  assign valid_396_reset = reset;
  assign valid_397_io_in = 1'h1;
  assign valid_397_io_enable = 1'h0;
  assign valid_397_clock = clock;
  assign valid_397_reset = reset;
  assign valid_398_io_in = 1'h1;
  assign valid_398_io_enable = 1'h0;
  assign valid_398_clock = clock;
  assign valid_398_reset = reset;
  assign valid_399_io_in = 1'h1;
  assign valid_399_io_enable = 1'h0;
  assign valid_399_clock = clock;
  assign valid_399_reset = reset;
  assign valid_400_io_in = 1'h1;
  assign valid_400_io_enable = 1'h0;
  assign valid_400_clock = clock;
  assign valid_400_reset = reset;
  assign valid_401_io_in = 1'h1;
  assign valid_401_io_enable = 1'h0;
  assign valid_401_clock = clock;
  assign valid_401_reset = reset;
  assign valid_402_io_in = 1'h1;
  assign valid_402_io_enable = 1'h0;
  assign valid_402_clock = clock;
  assign valid_402_reset = reset;
  assign valid_403_io_in = 1'h1;
  assign valid_403_io_enable = 1'h0;
  assign valid_403_clock = clock;
  assign valid_403_reset = reset;
  assign valid_404_io_in = 1'h1;
  assign valid_404_io_enable = 1'h0;
  assign valid_404_clock = clock;
  assign valid_404_reset = reset;
  assign valid_405_io_in = 1'h1;
  assign valid_405_io_enable = 1'h0;
  assign valid_405_clock = clock;
  assign valid_405_reset = reset;
  assign valid_406_io_in = 1'h1;
  assign valid_406_io_enable = 1'h0;
  assign valid_406_clock = clock;
  assign valid_406_reset = reset;
  assign valid_407_io_in = 1'h1;
  assign valid_407_io_enable = 1'h0;
  assign valid_407_clock = clock;
  assign valid_407_reset = reset;
  assign valid_408_io_in = 1'h1;
  assign valid_408_io_enable = 1'h0;
  assign valid_408_clock = clock;
  assign valid_408_reset = reset;
  assign valid_409_io_in = 1'h1;
  assign valid_409_io_enable = 1'h0;
  assign valid_409_clock = clock;
  assign valid_409_reset = reset;
  assign valid_410_io_in = 1'h1;
  assign valid_410_io_enable = 1'h0;
  assign valid_410_clock = clock;
  assign valid_410_reset = reset;
  assign valid_411_io_in = 1'h1;
  assign valid_411_io_enable = 1'h0;
  assign valid_411_clock = clock;
  assign valid_411_reset = reset;
  assign valid_412_io_in = 1'h1;
  assign valid_412_io_enable = 1'h0;
  assign valid_412_clock = clock;
  assign valid_412_reset = reset;
  assign valid_413_io_in = 1'h1;
  assign valid_413_io_enable = 1'h0;
  assign valid_413_clock = clock;
  assign valid_413_reset = reset;
  assign valid_414_io_in = 1'h1;
  assign valid_414_io_enable = 1'h0;
  assign valid_414_clock = clock;
  assign valid_414_reset = reset;
  assign valid_415_io_in = 1'h1;
  assign valid_415_io_enable = 1'h0;
  assign valid_415_clock = clock;
  assign valid_415_reset = reset;
  assign valid_416_io_in = 1'h1;
  assign valid_416_io_enable = 1'h0;
  assign valid_416_clock = clock;
  assign valid_416_reset = reset;
  assign valid_417_io_in = 1'h1;
  assign valid_417_io_enable = 1'h0;
  assign valid_417_clock = clock;
  assign valid_417_reset = reset;
  assign valid_418_io_in = 1'h1;
  assign valid_418_io_enable = 1'h0;
  assign valid_418_clock = clock;
  assign valid_418_reset = reset;
  assign valid_419_io_in = 1'h1;
  assign valid_419_io_enable = 1'h0;
  assign valid_419_clock = clock;
  assign valid_419_reset = reset;
  assign valid_420_io_in = 1'h1;
  assign valid_420_io_enable = 1'h0;
  assign valid_420_clock = clock;
  assign valid_420_reset = reset;
  assign valid_421_io_in = 1'h1;
  assign valid_421_io_enable = 1'h0;
  assign valid_421_clock = clock;
  assign valid_421_reset = reset;
  assign valid_422_io_in = 1'h1;
  assign valid_422_io_enable = 1'h0;
  assign valid_422_clock = clock;
  assign valid_422_reset = reset;
  assign valid_423_io_in = 1'h1;
  assign valid_423_io_enable = 1'h0;
  assign valid_423_clock = clock;
  assign valid_423_reset = reset;
  assign valid_424_io_in = 1'h1;
  assign valid_424_io_enable = 1'h0;
  assign valid_424_clock = clock;
  assign valid_424_reset = reset;
  assign valid_425_io_in = 1'h1;
  assign valid_425_io_enable = 1'h0;
  assign valid_425_clock = clock;
  assign valid_425_reset = reset;
  assign valid_426_io_in = 1'h1;
  assign valid_426_io_enable = 1'h0;
  assign valid_426_clock = clock;
  assign valid_426_reset = reset;
  assign valid_427_io_in = 1'h1;
  assign valid_427_io_enable = 1'h0;
  assign valid_427_clock = clock;
  assign valid_427_reset = reset;
  assign valid_428_io_in = 1'h1;
  assign valid_428_io_enable = 1'h0;
  assign valid_428_clock = clock;
  assign valid_428_reset = reset;
  assign valid_429_io_in = 1'h1;
  assign valid_429_io_enable = 1'h0;
  assign valid_429_clock = clock;
  assign valid_429_reset = reset;
  assign valid_430_io_in = 1'h1;
  assign valid_430_io_enable = 1'h0;
  assign valid_430_clock = clock;
  assign valid_430_reset = reset;
  assign valid_431_io_in = 1'h1;
  assign valid_431_io_enable = 1'h0;
  assign valid_431_clock = clock;
  assign valid_431_reset = reset;
  assign valid_432_io_in = 1'h1;
  assign valid_432_io_enable = 1'h0;
  assign valid_432_clock = clock;
  assign valid_432_reset = reset;
  assign valid_433_io_in = 1'h1;
  assign valid_433_io_enable = 1'h0;
  assign valid_433_clock = clock;
  assign valid_433_reset = reset;
  assign valid_434_io_in = 1'h1;
  assign valid_434_io_enable = 1'h0;
  assign valid_434_clock = clock;
  assign valid_434_reset = reset;
  assign valid_435_io_in = 1'h1;
  assign valid_435_io_enable = 1'h0;
  assign valid_435_clock = clock;
  assign valid_435_reset = reset;
  assign valid_436_io_in = 1'h1;
  assign valid_436_io_enable = 1'h0;
  assign valid_436_clock = clock;
  assign valid_436_reset = reset;
  assign valid_437_io_in = 1'h1;
  assign valid_437_io_enable = 1'h0;
  assign valid_437_clock = clock;
  assign valid_437_reset = reset;
  assign valid_438_io_in = 1'h1;
  assign valid_438_io_enable = 1'h0;
  assign valid_438_clock = clock;
  assign valid_438_reset = reset;
  assign valid_439_io_in = 1'h1;
  assign valid_439_io_enable = 1'h0;
  assign valid_439_clock = clock;
  assign valid_439_reset = reset;
  assign valid_440_io_in = 1'h1;
  assign valid_440_io_enable = 1'h0;
  assign valid_440_clock = clock;
  assign valid_440_reset = reset;
  assign valid_441_io_in = 1'h1;
  assign valid_441_io_enable = 1'h0;
  assign valid_441_clock = clock;
  assign valid_441_reset = reset;
  assign valid_442_io_in = 1'h1;
  assign valid_442_io_enable = 1'h0;
  assign valid_442_clock = clock;
  assign valid_442_reset = reset;
  assign valid_443_io_in = 1'h1;
  assign valid_443_io_enable = 1'h0;
  assign valid_443_clock = clock;
  assign valid_443_reset = reset;
  assign valid_444_io_in = 1'h1;
  assign valid_444_io_enable = 1'h0;
  assign valid_444_clock = clock;
  assign valid_444_reset = reset;
  assign valid_445_io_in = 1'h1;
  assign valid_445_io_enable = 1'h0;
  assign valid_445_clock = clock;
  assign valid_445_reset = reset;
  assign valid_446_io_in = 1'h1;
  assign valid_446_io_enable = 1'h0;
  assign valid_446_clock = clock;
  assign valid_446_reset = reset;
  assign valid_447_io_in = 1'h1;
  assign valid_447_io_enable = 1'h0;
  assign valid_447_clock = clock;
  assign valid_447_reset = reset;
  assign valid_448_io_in = 1'h1;
  assign valid_448_io_enable = 1'h0;
  assign valid_448_clock = clock;
  assign valid_448_reset = reset;
  assign valid_449_io_in = 1'h1;
  assign valid_449_io_enable = 1'h0;
  assign valid_449_clock = clock;
  assign valid_449_reset = reset;
  assign valid_450_io_in = 1'h1;
  assign valid_450_io_enable = 1'h0;
  assign valid_450_clock = clock;
  assign valid_450_reset = reset;
  assign valid_451_io_in = 1'h1;
  assign valid_451_io_enable = 1'h0;
  assign valid_451_clock = clock;
  assign valid_451_reset = reset;
  assign valid_452_io_in = 1'h1;
  assign valid_452_io_enable = 1'h0;
  assign valid_452_clock = clock;
  assign valid_452_reset = reset;
  assign valid_453_io_in = 1'h1;
  assign valid_453_io_enable = 1'h0;
  assign valid_453_clock = clock;
  assign valid_453_reset = reset;
  assign valid_454_io_in = 1'h1;
  assign valid_454_io_enable = 1'h0;
  assign valid_454_clock = clock;
  assign valid_454_reset = reset;
  assign valid_455_io_in = 1'h1;
  assign valid_455_io_enable = 1'h0;
  assign valid_455_clock = clock;
  assign valid_455_reset = reset;
  assign valid_456_io_in = 1'h1;
  assign valid_456_io_enable = 1'h0;
  assign valid_456_clock = clock;
  assign valid_456_reset = reset;
  assign valid_457_io_in = 1'h1;
  assign valid_457_io_enable = 1'h0;
  assign valid_457_clock = clock;
  assign valid_457_reset = reset;
  assign valid_458_io_in = 1'h1;
  assign valid_458_io_enable = 1'h0;
  assign valid_458_clock = clock;
  assign valid_458_reset = reset;
  assign valid_459_io_in = 1'h1;
  assign valid_459_io_enable = 1'h0;
  assign valid_459_clock = clock;
  assign valid_459_reset = reset;
  assign valid_460_io_in = 1'h1;
  assign valid_460_io_enable = 1'h0;
  assign valid_460_clock = clock;
  assign valid_460_reset = reset;
  assign valid_461_io_in = 1'h1;
  assign valid_461_io_enable = 1'h0;
  assign valid_461_clock = clock;
  assign valid_461_reset = reset;
  assign valid_462_io_in = 1'h1;
  assign valid_462_io_enable = 1'h0;
  assign valid_462_clock = clock;
  assign valid_462_reset = reset;
  assign valid_463_io_in = 1'h1;
  assign valid_463_io_enable = 1'h0;
  assign valid_463_clock = clock;
  assign valid_463_reset = reset;
  assign valid_464_io_in = 1'h1;
  assign valid_464_io_enable = 1'h0;
  assign valid_464_clock = clock;
  assign valid_464_reset = reset;
  assign valid_465_io_in = 1'h1;
  assign valid_465_io_enable = 1'h0;
  assign valid_465_clock = clock;
  assign valid_465_reset = reset;
  assign valid_466_io_in = 1'h1;
  assign valid_466_io_enable = 1'h0;
  assign valid_466_clock = clock;
  assign valid_466_reset = reset;
  assign valid_467_io_in = 1'h1;
  assign valid_467_io_enable = 1'h0;
  assign valid_467_clock = clock;
  assign valid_467_reset = reset;
  assign valid_468_io_in = 1'h1;
  assign valid_468_io_enable = 1'h0;
  assign valid_468_clock = clock;
  assign valid_468_reset = reset;
  assign valid_469_io_in = 1'h1;
  assign valid_469_io_enable = 1'h0;
  assign valid_469_clock = clock;
  assign valid_469_reset = reset;
  assign valid_470_io_in = 1'h1;
  assign valid_470_io_enable = 1'h0;
  assign valid_470_clock = clock;
  assign valid_470_reset = reset;
  assign valid_471_io_in = 1'h1;
  assign valid_471_io_enable = 1'h0;
  assign valid_471_clock = clock;
  assign valid_471_reset = reset;
  assign valid_472_io_in = 1'h1;
  assign valid_472_io_enable = 1'h0;
  assign valid_472_clock = clock;
  assign valid_472_reset = reset;
  assign valid_473_io_in = 1'h1;
  assign valid_473_io_enable = 1'h0;
  assign valid_473_clock = clock;
  assign valid_473_reset = reset;
  assign valid_474_io_in = 1'h1;
  assign valid_474_io_enable = 1'h0;
  assign valid_474_clock = clock;
  assign valid_474_reset = reset;
  assign valid_475_io_in = 1'h1;
  assign valid_475_io_enable = 1'h0;
  assign valid_475_clock = clock;
  assign valid_475_reset = reset;
  assign valid_476_io_in = 1'h1;
  assign valid_476_io_enable = 1'h0;
  assign valid_476_clock = clock;
  assign valid_476_reset = reset;
  assign valid_477_io_in = 1'h1;
  assign valid_477_io_enable = 1'h0;
  assign valid_477_clock = clock;
  assign valid_477_reset = reset;
  assign valid_478_io_in = 1'h1;
  assign valid_478_io_enable = 1'h0;
  assign valid_478_clock = clock;
  assign valid_478_reset = reset;
  assign valid_479_io_in = 1'h1;
  assign valid_479_io_enable = 1'h0;
  assign valid_479_clock = clock;
  assign valid_479_reset = reset;
  assign valid_480_io_in = 1'h1;
  assign valid_480_io_enable = 1'h0;
  assign valid_480_clock = clock;
  assign valid_480_reset = reset;
  assign valid_481_io_in = 1'h1;
  assign valid_481_io_enable = 1'h0;
  assign valid_481_clock = clock;
  assign valid_481_reset = reset;
  assign valid_482_io_in = 1'h1;
  assign valid_482_io_enable = 1'h0;
  assign valid_482_clock = clock;
  assign valid_482_reset = reset;
  assign valid_483_io_in = 1'h1;
  assign valid_483_io_enable = 1'h0;
  assign valid_483_clock = clock;
  assign valid_483_reset = reset;
  assign valid_484_io_in = 1'h1;
  assign valid_484_io_enable = 1'h0;
  assign valid_484_clock = clock;
  assign valid_484_reset = reset;
  assign valid_485_io_in = 1'h1;
  assign valid_485_io_enable = 1'h0;
  assign valid_485_clock = clock;
  assign valid_485_reset = reset;
  assign valid_486_io_in = 1'h1;
  assign valid_486_io_enable = 1'h0;
  assign valid_486_clock = clock;
  assign valid_486_reset = reset;
  assign valid_487_io_in = 1'h1;
  assign valid_487_io_enable = 1'h0;
  assign valid_487_clock = clock;
  assign valid_487_reset = reset;
  assign valid_488_io_in = 1'h1;
  assign valid_488_io_enable = 1'h0;
  assign valid_488_clock = clock;
  assign valid_488_reset = reset;
  assign valid_489_io_in = 1'h1;
  assign valid_489_io_enable = 1'h0;
  assign valid_489_clock = clock;
  assign valid_489_reset = reset;
  assign valid_490_io_in = 1'h1;
  assign valid_490_io_enable = 1'h0;
  assign valid_490_clock = clock;
  assign valid_490_reset = reset;
  assign valid_491_io_in = 1'h1;
  assign valid_491_io_enable = 1'h0;
  assign valid_491_clock = clock;
  assign valid_491_reset = reset;
  assign valid_492_io_in = 1'h1;
  assign valid_492_io_enable = 1'h0;
  assign valid_492_clock = clock;
  assign valid_492_reset = reset;
  assign valid_493_io_in = 1'h1;
  assign valid_493_io_enable = 1'h0;
  assign valid_493_clock = clock;
  assign valid_493_reset = reset;
  assign valid_494_io_in = 1'h1;
  assign valid_494_io_enable = 1'h0;
  assign valid_494_clock = clock;
  assign valid_494_reset = reset;
  assign valid_495_io_in = 1'h1;
  assign valid_495_io_enable = 1'h0;
  assign valid_495_clock = clock;
  assign valid_495_reset = reset;
  assign valid_496_io_in = 1'h1;
  assign valid_496_io_enable = 1'h0;
  assign valid_496_clock = clock;
  assign valid_496_reset = reset;
  assign valid_497_io_in = 1'h1;
  assign valid_497_io_enable = 1'h0;
  assign valid_497_clock = clock;
  assign valid_497_reset = reset;
  assign valid_498_io_in = 1'h1;
  assign valid_498_io_enable = 1'h0;
  assign valid_498_clock = clock;
  assign valid_498_reset = reset;
  assign valid_499_io_in = 1'h1;
  assign valid_499_io_enable = 1'h0;
  assign valid_499_clock = clock;
  assign valid_499_reset = reset;
  assign valid_500_io_in = 1'h1;
  assign valid_500_io_enable = 1'h0;
  assign valid_500_clock = clock;
  assign valid_500_reset = reset;
  assign valid_501_io_in = 1'h1;
  assign valid_501_io_enable = 1'h0;
  assign valid_501_clock = clock;
  assign valid_501_reset = reset;
  assign valid_502_io_in = 1'h1;
  assign valid_502_io_enable = 1'h0;
  assign valid_502_clock = clock;
  assign valid_502_reset = reset;
  assign valid_503_io_in = 1'h1;
  assign valid_503_io_enable = 1'h0;
  assign valid_503_clock = clock;
  assign valid_503_reset = reset;
  assign valid_504_io_in = 1'h1;
  assign valid_504_io_enable = 1'h0;
  assign valid_504_clock = clock;
  assign valid_504_reset = reset;
  assign valid_505_io_in = 1'h1;
  assign valid_505_io_enable = 1'h0;
  assign valid_505_clock = clock;
  assign valid_505_reset = reset;
  assign valid_506_io_in = 1'h1;
  assign valid_506_io_enable = 1'h0;
  assign valid_506_clock = clock;
  assign valid_506_reset = reset;
  assign valid_507_io_in = 1'h1;
  assign valid_507_io_enable = 1'h0;
  assign valid_507_clock = clock;
  assign valid_507_reset = reset;
  assign valid_508_io_in = 1'h1;
  assign valid_508_io_enable = 1'h0;
  assign valid_508_clock = clock;
  assign valid_508_reset = reset;
  assign valid_509_io_in = 1'h1;
  assign valid_509_io_enable = 1'h0;
  assign valid_509_clock = clock;
  assign valid_509_reset = reset;
  assign valid_510_io_in = 1'h1;
  assign valid_510_io_enable = 1'h0;
  assign valid_510_clock = clock;
  assign valid_510_reset = reset;
  assign valid_511_io_in = 1'h1;
  assign valid_511_io_enable = 1'h0;
  assign valid_511_clock = clock;
  assign valid_511_reset = reset;
  assign tags_0_clock = clock;
  assign tags_0_reset = reset;
  assign tags_1_clock = clock;
  assign tags_1_reset = reset;
  assign tags_2_clock = clock;
  assign tags_2_reset = reset;
  assign tags_3_clock = clock;
  assign tags_3_reset = reset;
  assign tags_4_clock = clock;
  assign tags_4_reset = reset;
  assign tags_5_clock = clock;
  assign tags_5_reset = reset;
  assign tags_6_clock = clock;
  assign tags_6_reset = reset;
  assign tags_7_clock = clock;
  assign tags_7_reset = reset;
  assign tags_8_clock = clock;
  assign tags_8_reset = reset;
  assign tags_9_clock = clock;
  assign tags_9_reset = reset;
  assign tags_10_clock = clock;
  assign tags_10_reset = reset;
  assign tags_11_clock = clock;
  assign tags_11_reset = reset;
  assign tags_12_clock = clock;
  assign tags_12_reset = reset;
  assign tags_13_clock = clock;
  assign tags_13_reset = reset;
  assign tags_14_clock = clock;
  assign tags_14_reset = reset;
  assign tags_15_clock = clock;
  assign tags_15_reset = reset;
  assign tags_16_clock = clock;
  assign tags_16_reset = reset;
  assign tags_17_clock = clock;
  assign tags_17_reset = reset;
  assign tags_18_clock = clock;
  assign tags_18_reset = reset;
  assign tags_19_clock = clock;
  assign tags_19_reset = reset;
  assign tags_20_clock = clock;
  assign tags_20_reset = reset;
  assign tags_21_clock = clock;
  assign tags_21_reset = reset;
  assign tags_22_clock = clock;
  assign tags_22_reset = reset;
  assign tags_23_clock = clock;
  assign tags_23_reset = reset;
  assign tags_24_clock = clock;
  assign tags_24_reset = reset;
  assign tags_25_clock = clock;
  assign tags_25_reset = reset;
  assign tags_26_clock = clock;
  assign tags_26_reset = reset;
  assign tags_27_clock = clock;
  assign tags_27_reset = reset;
  assign tags_28_clock = clock;
  assign tags_28_reset = reset;
  assign tags_29_clock = clock;
  assign tags_29_reset = reset;
  assign tags_30_clock = clock;
  assign tags_30_reset = reset;
  assign tags_31_clock = clock;
  assign tags_31_reset = reset;
  assign tags_32_clock = clock;
  assign tags_32_reset = reset;
  assign tags_33_clock = clock;
  assign tags_33_reset = reset;
  assign tags_34_clock = clock;
  assign tags_34_reset = reset;
  assign tags_35_clock = clock;
  assign tags_35_reset = reset;
  assign tags_36_clock = clock;
  assign tags_36_reset = reset;
  assign tags_37_clock = clock;
  assign tags_37_reset = reset;
  assign tags_38_clock = clock;
  assign tags_38_reset = reset;
  assign tags_39_clock = clock;
  assign tags_39_reset = reset;
  assign tags_40_clock = clock;
  assign tags_40_reset = reset;
  assign tags_41_clock = clock;
  assign tags_41_reset = reset;
  assign tags_42_clock = clock;
  assign tags_42_reset = reset;
  assign tags_43_clock = clock;
  assign tags_43_reset = reset;
  assign tags_44_clock = clock;
  assign tags_44_reset = reset;
  assign tags_45_clock = clock;
  assign tags_45_reset = reset;
  assign tags_46_clock = clock;
  assign tags_46_reset = reset;
  assign tags_47_clock = clock;
  assign tags_47_reset = reset;
  assign tags_48_clock = clock;
  assign tags_48_reset = reset;
  assign tags_49_clock = clock;
  assign tags_49_reset = reset;
  assign tags_50_clock = clock;
  assign tags_50_reset = reset;
  assign tags_51_clock = clock;
  assign tags_51_reset = reset;
  assign tags_52_clock = clock;
  assign tags_52_reset = reset;
  assign tags_53_clock = clock;
  assign tags_53_reset = reset;
  assign tags_54_clock = clock;
  assign tags_54_reset = reset;
  assign tags_55_clock = clock;
  assign tags_55_reset = reset;
  assign tags_56_clock = clock;
  assign tags_56_reset = reset;
  assign tags_57_clock = clock;
  assign tags_57_reset = reset;
  assign tags_58_clock = clock;
  assign tags_58_reset = reset;
  assign tags_59_clock = clock;
  assign tags_59_reset = reset;
  assign tags_60_clock = clock;
  assign tags_60_reset = reset;
  assign tags_61_clock = clock;
  assign tags_61_reset = reset;
  assign tags_62_clock = clock;
  assign tags_62_reset = reset;
  assign tags_63_clock = clock;
  assign tags_63_reset = reset;
  assign tags_64_clock = clock;
  assign tags_64_reset = reset;
  assign tags_65_clock = clock;
  assign tags_65_reset = reset;
  assign tags_66_clock = clock;
  assign tags_66_reset = reset;
  assign tags_67_clock = clock;
  assign tags_67_reset = reset;
  assign tags_68_clock = clock;
  assign tags_68_reset = reset;
  assign tags_69_clock = clock;
  assign tags_69_reset = reset;
  assign tags_70_clock = clock;
  assign tags_70_reset = reset;
  assign tags_71_clock = clock;
  assign tags_71_reset = reset;
  assign tags_72_clock = clock;
  assign tags_72_reset = reset;
  assign tags_73_clock = clock;
  assign tags_73_reset = reset;
  assign tags_74_clock = clock;
  assign tags_74_reset = reset;
  assign tags_75_clock = clock;
  assign tags_75_reset = reset;
  assign tags_76_clock = clock;
  assign tags_76_reset = reset;
  assign tags_77_clock = clock;
  assign tags_77_reset = reset;
  assign tags_78_clock = clock;
  assign tags_78_reset = reset;
  assign tags_79_clock = clock;
  assign tags_79_reset = reset;
  assign tags_80_clock = clock;
  assign tags_80_reset = reset;
  assign tags_81_clock = clock;
  assign tags_81_reset = reset;
  assign tags_82_clock = clock;
  assign tags_82_reset = reset;
  assign tags_83_clock = clock;
  assign tags_83_reset = reset;
  assign tags_84_clock = clock;
  assign tags_84_reset = reset;
  assign tags_85_clock = clock;
  assign tags_85_reset = reset;
  assign tags_86_clock = clock;
  assign tags_86_reset = reset;
  assign tags_87_clock = clock;
  assign tags_87_reset = reset;
  assign tags_88_clock = clock;
  assign tags_88_reset = reset;
  assign tags_89_clock = clock;
  assign tags_89_reset = reset;
  assign tags_90_clock = clock;
  assign tags_90_reset = reset;
  assign tags_91_clock = clock;
  assign tags_91_reset = reset;
  assign tags_92_clock = clock;
  assign tags_92_reset = reset;
  assign tags_93_clock = clock;
  assign tags_93_reset = reset;
  assign tags_94_clock = clock;
  assign tags_94_reset = reset;
  assign tags_95_clock = clock;
  assign tags_95_reset = reset;
  assign tags_96_clock = clock;
  assign tags_96_reset = reset;
  assign tags_97_clock = clock;
  assign tags_97_reset = reset;
  assign tags_98_clock = clock;
  assign tags_98_reset = reset;
  assign tags_99_clock = clock;
  assign tags_99_reset = reset;
  assign tags_100_clock = clock;
  assign tags_100_reset = reset;
  assign tags_101_clock = clock;
  assign tags_101_reset = reset;
  assign tags_102_clock = clock;
  assign tags_102_reset = reset;
  assign tags_103_clock = clock;
  assign tags_103_reset = reset;
  assign tags_104_clock = clock;
  assign tags_104_reset = reset;
  assign tags_105_clock = clock;
  assign tags_105_reset = reset;
  assign tags_106_clock = clock;
  assign tags_106_reset = reset;
  assign tags_107_clock = clock;
  assign tags_107_reset = reset;
  assign tags_108_clock = clock;
  assign tags_108_reset = reset;
  assign tags_109_clock = clock;
  assign tags_109_reset = reset;
  assign tags_110_clock = clock;
  assign tags_110_reset = reset;
  assign tags_111_clock = clock;
  assign tags_111_reset = reset;
  assign tags_112_clock = clock;
  assign tags_112_reset = reset;
  assign tags_113_clock = clock;
  assign tags_113_reset = reset;
  assign tags_114_clock = clock;
  assign tags_114_reset = reset;
  assign tags_115_clock = clock;
  assign tags_115_reset = reset;
  assign tags_116_clock = clock;
  assign tags_116_reset = reset;
  assign tags_117_clock = clock;
  assign tags_117_reset = reset;
  assign tags_118_clock = clock;
  assign tags_118_reset = reset;
  assign tags_119_clock = clock;
  assign tags_119_reset = reset;
  assign tags_120_clock = clock;
  assign tags_120_reset = reset;
  assign tags_121_clock = clock;
  assign tags_121_reset = reset;
  assign tags_122_clock = clock;
  assign tags_122_reset = reset;
  assign tags_123_clock = clock;
  assign tags_123_reset = reset;
  assign tags_124_clock = clock;
  assign tags_124_reset = reset;
  assign tags_125_clock = clock;
  assign tags_125_reset = reset;
  assign tags_126_clock = clock;
  assign tags_126_reset = reset;
  assign tags_127_clock = clock;
  assign tags_127_reset = reset;
  assign tags_128_clock = clock;
  assign tags_128_reset = reset;
  assign tags_129_clock = clock;
  assign tags_129_reset = reset;
  assign tags_130_clock = clock;
  assign tags_130_reset = reset;
  assign tags_131_clock = clock;
  assign tags_131_reset = reset;
  assign tags_132_clock = clock;
  assign tags_132_reset = reset;
  assign tags_133_clock = clock;
  assign tags_133_reset = reset;
  assign tags_134_clock = clock;
  assign tags_134_reset = reset;
  assign tags_135_clock = clock;
  assign tags_135_reset = reset;
  assign tags_136_clock = clock;
  assign tags_136_reset = reset;
  assign tags_137_clock = clock;
  assign tags_137_reset = reset;
  assign tags_138_clock = clock;
  assign tags_138_reset = reset;
  assign tags_139_clock = clock;
  assign tags_139_reset = reset;
  assign tags_140_clock = clock;
  assign tags_140_reset = reset;
  assign tags_141_clock = clock;
  assign tags_141_reset = reset;
  assign tags_142_clock = clock;
  assign tags_142_reset = reset;
  assign tags_143_clock = clock;
  assign tags_143_reset = reset;
  assign tags_144_clock = clock;
  assign tags_144_reset = reset;
  assign tags_145_clock = clock;
  assign tags_145_reset = reset;
  assign tags_146_clock = clock;
  assign tags_146_reset = reset;
  assign tags_147_clock = clock;
  assign tags_147_reset = reset;
  assign tags_148_clock = clock;
  assign tags_148_reset = reset;
  assign tags_149_clock = clock;
  assign tags_149_reset = reset;
  assign tags_150_clock = clock;
  assign tags_150_reset = reset;
  assign tags_151_clock = clock;
  assign tags_151_reset = reset;
  assign tags_152_clock = clock;
  assign tags_152_reset = reset;
  assign tags_153_clock = clock;
  assign tags_153_reset = reset;
  assign tags_154_clock = clock;
  assign tags_154_reset = reset;
  assign tags_155_clock = clock;
  assign tags_155_reset = reset;
  assign tags_156_clock = clock;
  assign tags_156_reset = reset;
  assign tags_157_clock = clock;
  assign tags_157_reset = reset;
  assign tags_158_clock = clock;
  assign tags_158_reset = reset;
  assign tags_159_clock = clock;
  assign tags_159_reset = reset;
  assign tags_160_clock = clock;
  assign tags_160_reset = reset;
  assign tags_161_clock = clock;
  assign tags_161_reset = reset;
  assign tags_162_clock = clock;
  assign tags_162_reset = reset;
  assign tags_163_clock = clock;
  assign tags_163_reset = reset;
  assign tags_164_clock = clock;
  assign tags_164_reset = reset;
  assign tags_165_clock = clock;
  assign tags_165_reset = reset;
  assign tags_166_clock = clock;
  assign tags_166_reset = reset;
  assign tags_167_clock = clock;
  assign tags_167_reset = reset;
  assign tags_168_clock = clock;
  assign tags_168_reset = reset;
  assign tags_169_clock = clock;
  assign tags_169_reset = reset;
  assign tags_170_clock = clock;
  assign tags_170_reset = reset;
  assign tags_171_clock = clock;
  assign tags_171_reset = reset;
  assign tags_172_clock = clock;
  assign tags_172_reset = reset;
  assign tags_173_clock = clock;
  assign tags_173_reset = reset;
  assign tags_174_clock = clock;
  assign tags_174_reset = reset;
  assign tags_175_clock = clock;
  assign tags_175_reset = reset;
  assign tags_176_clock = clock;
  assign tags_176_reset = reset;
  assign tags_177_clock = clock;
  assign tags_177_reset = reset;
  assign tags_178_clock = clock;
  assign tags_178_reset = reset;
  assign tags_179_clock = clock;
  assign tags_179_reset = reset;
  assign tags_180_clock = clock;
  assign tags_180_reset = reset;
  assign tags_181_clock = clock;
  assign tags_181_reset = reset;
  assign tags_182_clock = clock;
  assign tags_182_reset = reset;
  assign tags_183_clock = clock;
  assign tags_183_reset = reset;
  assign tags_184_clock = clock;
  assign tags_184_reset = reset;
  assign tags_185_clock = clock;
  assign tags_185_reset = reset;
  assign tags_186_clock = clock;
  assign tags_186_reset = reset;
  assign tags_187_clock = clock;
  assign tags_187_reset = reset;
  assign tags_188_clock = clock;
  assign tags_188_reset = reset;
  assign tags_189_clock = clock;
  assign tags_189_reset = reset;
  assign tags_190_clock = clock;
  assign tags_190_reset = reset;
  assign tags_191_clock = clock;
  assign tags_191_reset = reset;
  assign tags_192_clock = clock;
  assign tags_192_reset = reset;
  assign tags_193_clock = clock;
  assign tags_193_reset = reset;
  assign tags_194_clock = clock;
  assign tags_194_reset = reset;
  assign tags_195_clock = clock;
  assign tags_195_reset = reset;
  assign tags_196_clock = clock;
  assign tags_196_reset = reset;
  assign tags_197_clock = clock;
  assign tags_197_reset = reset;
  assign tags_198_clock = clock;
  assign tags_198_reset = reset;
  assign tags_199_clock = clock;
  assign tags_199_reset = reset;
  assign tags_200_clock = clock;
  assign tags_200_reset = reset;
  assign tags_201_clock = clock;
  assign tags_201_reset = reset;
  assign tags_202_clock = clock;
  assign tags_202_reset = reset;
  assign tags_203_clock = clock;
  assign tags_203_reset = reset;
  assign tags_204_clock = clock;
  assign tags_204_reset = reset;
  assign tags_205_clock = clock;
  assign tags_205_reset = reset;
  assign tags_206_clock = clock;
  assign tags_206_reset = reset;
  assign tags_207_clock = clock;
  assign tags_207_reset = reset;
  assign tags_208_clock = clock;
  assign tags_208_reset = reset;
  assign tags_209_clock = clock;
  assign tags_209_reset = reset;
  assign tags_210_clock = clock;
  assign tags_210_reset = reset;
  assign tags_211_clock = clock;
  assign tags_211_reset = reset;
  assign tags_212_clock = clock;
  assign tags_212_reset = reset;
  assign tags_213_clock = clock;
  assign tags_213_reset = reset;
  assign tags_214_clock = clock;
  assign tags_214_reset = reset;
  assign tags_215_clock = clock;
  assign tags_215_reset = reset;
  assign tags_216_clock = clock;
  assign tags_216_reset = reset;
  assign tags_217_clock = clock;
  assign tags_217_reset = reset;
  assign tags_218_clock = clock;
  assign tags_218_reset = reset;
  assign tags_219_clock = clock;
  assign tags_219_reset = reset;
  assign tags_220_clock = clock;
  assign tags_220_reset = reset;
  assign tags_221_clock = clock;
  assign tags_221_reset = reset;
  assign tags_222_clock = clock;
  assign tags_222_reset = reset;
  assign tags_223_clock = clock;
  assign tags_223_reset = reset;
  assign tags_224_clock = clock;
  assign tags_224_reset = reset;
  assign tags_225_clock = clock;
  assign tags_225_reset = reset;
  assign tags_226_clock = clock;
  assign tags_226_reset = reset;
  assign tags_227_clock = clock;
  assign tags_227_reset = reset;
  assign tags_228_clock = clock;
  assign tags_228_reset = reset;
  assign tags_229_clock = clock;
  assign tags_229_reset = reset;
  assign tags_230_clock = clock;
  assign tags_230_reset = reset;
  assign tags_231_clock = clock;
  assign tags_231_reset = reset;
  assign tags_232_clock = clock;
  assign tags_232_reset = reset;
  assign tags_233_clock = clock;
  assign tags_233_reset = reset;
  assign tags_234_clock = clock;
  assign tags_234_reset = reset;
  assign tags_235_clock = clock;
  assign tags_235_reset = reset;
  assign tags_236_clock = clock;
  assign tags_236_reset = reset;
  assign tags_237_clock = clock;
  assign tags_237_reset = reset;
  assign tags_238_clock = clock;
  assign tags_238_reset = reset;
  assign tags_239_clock = clock;
  assign tags_239_reset = reset;
  assign tags_240_clock = clock;
  assign tags_240_reset = reset;
  assign tags_241_clock = clock;
  assign tags_241_reset = reset;
  assign tags_242_clock = clock;
  assign tags_242_reset = reset;
  assign tags_243_clock = clock;
  assign tags_243_reset = reset;
  assign tags_244_clock = clock;
  assign tags_244_reset = reset;
  assign tags_245_clock = clock;
  assign tags_245_reset = reset;
  assign tags_246_clock = clock;
  assign tags_246_reset = reset;
  assign tags_247_clock = clock;
  assign tags_247_reset = reset;
  assign tags_248_clock = clock;
  assign tags_248_reset = reset;
  assign tags_249_clock = clock;
  assign tags_249_reset = reset;
  assign tags_250_clock = clock;
  assign tags_250_reset = reset;
  assign tags_251_clock = clock;
  assign tags_251_reset = reset;
  assign tags_252_clock = clock;
  assign tags_252_reset = reset;
  assign tags_253_clock = clock;
  assign tags_253_reset = reset;
  assign tags_254_clock = clock;
  assign tags_254_reset = reset;
  assign tags_255_clock = clock;
  assign tags_255_reset = reset;
  assign tags_256_clock = clock;
  assign tags_256_reset = reset;
  assign tags_257_clock = clock;
  assign tags_257_reset = reset;
  assign tags_258_clock = clock;
  assign tags_258_reset = reset;
  assign tags_259_clock = clock;
  assign tags_259_reset = reset;
  assign tags_260_clock = clock;
  assign tags_260_reset = reset;
  assign tags_261_clock = clock;
  assign tags_261_reset = reset;
  assign tags_262_clock = clock;
  assign tags_262_reset = reset;
  assign tags_263_clock = clock;
  assign tags_263_reset = reset;
  assign tags_264_clock = clock;
  assign tags_264_reset = reset;
  assign tags_265_clock = clock;
  assign tags_265_reset = reset;
  assign tags_266_clock = clock;
  assign tags_266_reset = reset;
  assign tags_267_clock = clock;
  assign tags_267_reset = reset;
  assign tags_268_clock = clock;
  assign tags_268_reset = reset;
  assign tags_269_clock = clock;
  assign tags_269_reset = reset;
  assign tags_270_clock = clock;
  assign tags_270_reset = reset;
  assign tags_271_clock = clock;
  assign tags_271_reset = reset;
  assign tags_272_clock = clock;
  assign tags_272_reset = reset;
  assign tags_273_clock = clock;
  assign tags_273_reset = reset;
  assign tags_274_clock = clock;
  assign tags_274_reset = reset;
  assign tags_275_clock = clock;
  assign tags_275_reset = reset;
  assign tags_276_clock = clock;
  assign tags_276_reset = reset;
  assign tags_277_clock = clock;
  assign tags_277_reset = reset;
  assign tags_278_clock = clock;
  assign tags_278_reset = reset;
  assign tags_279_clock = clock;
  assign tags_279_reset = reset;
  assign tags_280_clock = clock;
  assign tags_280_reset = reset;
  assign tags_281_clock = clock;
  assign tags_281_reset = reset;
  assign tags_282_clock = clock;
  assign tags_282_reset = reset;
  assign tags_283_clock = clock;
  assign tags_283_reset = reset;
  assign tags_284_clock = clock;
  assign tags_284_reset = reset;
  assign tags_285_clock = clock;
  assign tags_285_reset = reset;
  assign tags_286_clock = clock;
  assign tags_286_reset = reset;
  assign tags_287_clock = clock;
  assign tags_287_reset = reset;
  assign tags_288_clock = clock;
  assign tags_288_reset = reset;
  assign tags_289_clock = clock;
  assign tags_289_reset = reset;
  assign tags_290_clock = clock;
  assign tags_290_reset = reset;
  assign tags_291_clock = clock;
  assign tags_291_reset = reset;
  assign tags_292_clock = clock;
  assign tags_292_reset = reset;
  assign tags_293_clock = clock;
  assign tags_293_reset = reset;
  assign tags_294_clock = clock;
  assign tags_294_reset = reset;
  assign tags_295_clock = clock;
  assign tags_295_reset = reset;
  assign tags_296_clock = clock;
  assign tags_296_reset = reset;
  assign tags_297_clock = clock;
  assign tags_297_reset = reset;
  assign tags_298_clock = clock;
  assign tags_298_reset = reset;
  assign tags_299_clock = clock;
  assign tags_299_reset = reset;
  assign tags_300_clock = clock;
  assign tags_300_reset = reset;
  assign tags_301_clock = clock;
  assign tags_301_reset = reset;
  assign tags_302_clock = clock;
  assign tags_302_reset = reset;
  assign tags_303_clock = clock;
  assign tags_303_reset = reset;
  assign tags_304_clock = clock;
  assign tags_304_reset = reset;
  assign tags_305_clock = clock;
  assign tags_305_reset = reset;
  assign tags_306_clock = clock;
  assign tags_306_reset = reset;
  assign tags_307_clock = clock;
  assign tags_307_reset = reset;
  assign tags_308_clock = clock;
  assign tags_308_reset = reset;
  assign tags_309_clock = clock;
  assign tags_309_reset = reset;
  assign tags_310_clock = clock;
  assign tags_310_reset = reset;
  assign tags_311_clock = clock;
  assign tags_311_reset = reset;
  assign tags_312_clock = clock;
  assign tags_312_reset = reset;
  assign tags_313_clock = clock;
  assign tags_313_reset = reset;
  assign tags_314_clock = clock;
  assign tags_314_reset = reset;
  assign tags_315_clock = clock;
  assign tags_315_reset = reset;
  assign tags_316_clock = clock;
  assign tags_316_reset = reset;
  assign tags_317_clock = clock;
  assign tags_317_reset = reset;
  assign tags_318_clock = clock;
  assign tags_318_reset = reset;
  assign tags_319_clock = clock;
  assign tags_319_reset = reset;
  assign tags_320_clock = clock;
  assign tags_320_reset = reset;
  assign tags_321_clock = clock;
  assign tags_321_reset = reset;
  assign tags_322_clock = clock;
  assign tags_322_reset = reset;
  assign tags_323_clock = clock;
  assign tags_323_reset = reset;
  assign tags_324_clock = clock;
  assign tags_324_reset = reset;
  assign tags_325_clock = clock;
  assign tags_325_reset = reset;
  assign tags_326_clock = clock;
  assign tags_326_reset = reset;
  assign tags_327_clock = clock;
  assign tags_327_reset = reset;
  assign tags_328_clock = clock;
  assign tags_328_reset = reset;
  assign tags_329_clock = clock;
  assign tags_329_reset = reset;
  assign tags_330_clock = clock;
  assign tags_330_reset = reset;
  assign tags_331_clock = clock;
  assign tags_331_reset = reset;
  assign tags_332_clock = clock;
  assign tags_332_reset = reset;
  assign tags_333_clock = clock;
  assign tags_333_reset = reset;
  assign tags_334_clock = clock;
  assign tags_334_reset = reset;
  assign tags_335_clock = clock;
  assign tags_335_reset = reset;
  assign tags_336_clock = clock;
  assign tags_336_reset = reset;
  assign tags_337_clock = clock;
  assign tags_337_reset = reset;
  assign tags_338_clock = clock;
  assign tags_338_reset = reset;
  assign tags_339_clock = clock;
  assign tags_339_reset = reset;
  assign tags_340_clock = clock;
  assign tags_340_reset = reset;
  assign tags_341_clock = clock;
  assign tags_341_reset = reset;
  assign tags_342_clock = clock;
  assign tags_342_reset = reset;
  assign tags_343_clock = clock;
  assign tags_343_reset = reset;
  assign tags_344_clock = clock;
  assign tags_344_reset = reset;
  assign tags_345_clock = clock;
  assign tags_345_reset = reset;
  assign tags_346_clock = clock;
  assign tags_346_reset = reset;
  assign tags_347_clock = clock;
  assign tags_347_reset = reset;
  assign tags_348_clock = clock;
  assign tags_348_reset = reset;
  assign tags_349_clock = clock;
  assign tags_349_reset = reset;
  assign tags_350_clock = clock;
  assign tags_350_reset = reset;
  assign tags_351_clock = clock;
  assign tags_351_reset = reset;
  assign tags_352_clock = clock;
  assign tags_352_reset = reset;
  assign tags_353_clock = clock;
  assign tags_353_reset = reset;
  assign tags_354_clock = clock;
  assign tags_354_reset = reset;
  assign tags_355_clock = clock;
  assign tags_355_reset = reset;
  assign tags_356_clock = clock;
  assign tags_356_reset = reset;
  assign tags_357_clock = clock;
  assign tags_357_reset = reset;
  assign tags_358_clock = clock;
  assign tags_358_reset = reset;
  assign tags_359_clock = clock;
  assign tags_359_reset = reset;
  assign tags_360_clock = clock;
  assign tags_360_reset = reset;
  assign tags_361_clock = clock;
  assign tags_361_reset = reset;
  assign tags_362_clock = clock;
  assign tags_362_reset = reset;
  assign tags_363_clock = clock;
  assign tags_363_reset = reset;
  assign tags_364_clock = clock;
  assign tags_364_reset = reset;
  assign tags_365_clock = clock;
  assign tags_365_reset = reset;
  assign tags_366_clock = clock;
  assign tags_366_reset = reset;
  assign tags_367_clock = clock;
  assign tags_367_reset = reset;
  assign tags_368_clock = clock;
  assign tags_368_reset = reset;
  assign tags_369_clock = clock;
  assign tags_369_reset = reset;
  assign tags_370_clock = clock;
  assign tags_370_reset = reset;
  assign tags_371_clock = clock;
  assign tags_371_reset = reset;
  assign tags_372_clock = clock;
  assign tags_372_reset = reset;
  assign tags_373_clock = clock;
  assign tags_373_reset = reset;
  assign tags_374_clock = clock;
  assign tags_374_reset = reset;
  assign tags_375_clock = clock;
  assign tags_375_reset = reset;
  assign tags_376_clock = clock;
  assign tags_376_reset = reset;
  assign tags_377_clock = clock;
  assign tags_377_reset = reset;
  assign tags_378_clock = clock;
  assign tags_378_reset = reset;
  assign tags_379_clock = clock;
  assign tags_379_reset = reset;
  assign tags_380_clock = clock;
  assign tags_380_reset = reset;
  assign tags_381_clock = clock;
  assign tags_381_reset = reset;
  assign tags_382_clock = clock;
  assign tags_382_reset = reset;
  assign tags_383_clock = clock;
  assign tags_383_reset = reset;
  assign tags_384_clock = clock;
  assign tags_384_reset = reset;
  assign tags_385_clock = clock;
  assign tags_385_reset = reset;
  assign tags_386_clock = clock;
  assign tags_386_reset = reset;
  assign tags_387_clock = clock;
  assign tags_387_reset = reset;
  assign tags_388_clock = clock;
  assign tags_388_reset = reset;
  assign tags_389_clock = clock;
  assign tags_389_reset = reset;
  assign tags_390_clock = clock;
  assign tags_390_reset = reset;
  assign tags_391_clock = clock;
  assign tags_391_reset = reset;
  assign tags_392_clock = clock;
  assign tags_392_reset = reset;
  assign tags_393_clock = clock;
  assign tags_393_reset = reset;
  assign tags_394_clock = clock;
  assign tags_394_reset = reset;
  assign tags_395_clock = clock;
  assign tags_395_reset = reset;
  assign tags_396_clock = clock;
  assign tags_396_reset = reset;
  assign tags_397_clock = clock;
  assign tags_397_reset = reset;
  assign tags_398_clock = clock;
  assign tags_398_reset = reset;
  assign tags_399_clock = clock;
  assign tags_399_reset = reset;
  assign tags_400_clock = clock;
  assign tags_400_reset = reset;
  assign tags_401_clock = clock;
  assign tags_401_reset = reset;
  assign tags_402_clock = clock;
  assign tags_402_reset = reset;
  assign tags_403_clock = clock;
  assign tags_403_reset = reset;
  assign tags_404_clock = clock;
  assign tags_404_reset = reset;
  assign tags_405_clock = clock;
  assign tags_405_reset = reset;
  assign tags_406_clock = clock;
  assign tags_406_reset = reset;
  assign tags_407_clock = clock;
  assign tags_407_reset = reset;
  assign tags_408_clock = clock;
  assign tags_408_reset = reset;
  assign tags_409_clock = clock;
  assign tags_409_reset = reset;
  assign tags_410_clock = clock;
  assign tags_410_reset = reset;
  assign tags_411_clock = clock;
  assign tags_411_reset = reset;
  assign tags_412_clock = clock;
  assign tags_412_reset = reset;
  assign tags_413_clock = clock;
  assign tags_413_reset = reset;
  assign tags_414_clock = clock;
  assign tags_414_reset = reset;
  assign tags_415_clock = clock;
  assign tags_415_reset = reset;
  assign tags_416_clock = clock;
  assign tags_416_reset = reset;
  assign tags_417_clock = clock;
  assign tags_417_reset = reset;
  assign tags_418_clock = clock;
  assign tags_418_reset = reset;
  assign tags_419_clock = clock;
  assign tags_419_reset = reset;
  assign tags_420_clock = clock;
  assign tags_420_reset = reset;
  assign tags_421_clock = clock;
  assign tags_421_reset = reset;
  assign tags_422_clock = clock;
  assign tags_422_reset = reset;
  assign tags_423_clock = clock;
  assign tags_423_reset = reset;
  assign tags_424_clock = clock;
  assign tags_424_reset = reset;
  assign tags_425_clock = clock;
  assign tags_425_reset = reset;
  assign tags_426_clock = clock;
  assign tags_426_reset = reset;
  assign tags_427_clock = clock;
  assign tags_427_reset = reset;
  assign tags_428_clock = clock;
  assign tags_428_reset = reset;
  assign tags_429_clock = clock;
  assign tags_429_reset = reset;
  assign tags_430_clock = clock;
  assign tags_430_reset = reset;
  assign tags_431_clock = clock;
  assign tags_431_reset = reset;
  assign tags_432_clock = clock;
  assign tags_432_reset = reset;
  assign tags_433_clock = clock;
  assign tags_433_reset = reset;
  assign tags_434_clock = clock;
  assign tags_434_reset = reset;
  assign tags_435_clock = clock;
  assign tags_435_reset = reset;
  assign tags_436_clock = clock;
  assign tags_436_reset = reset;
  assign tags_437_clock = clock;
  assign tags_437_reset = reset;
  assign tags_438_clock = clock;
  assign tags_438_reset = reset;
  assign tags_439_clock = clock;
  assign tags_439_reset = reset;
  assign tags_440_clock = clock;
  assign tags_440_reset = reset;
  assign tags_441_clock = clock;
  assign tags_441_reset = reset;
  assign tags_442_clock = clock;
  assign tags_442_reset = reset;
  assign tags_443_clock = clock;
  assign tags_443_reset = reset;
  assign tags_444_clock = clock;
  assign tags_444_reset = reset;
  assign tags_445_clock = clock;
  assign tags_445_reset = reset;
  assign tags_446_clock = clock;
  assign tags_446_reset = reset;
  assign tags_447_clock = clock;
  assign tags_447_reset = reset;
  assign tags_448_clock = clock;
  assign tags_448_reset = reset;
  assign tags_449_clock = clock;
  assign tags_449_reset = reset;
  assign tags_450_clock = clock;
  assign tags_450_reset = reset;
  assign tags_451_clock = clock;
  assign tags_451_reset = reset;
  assign tags_452_clock = clock;
  assign tags_452_reset = reset;
  assign tags_453_clock = clock;
  assign tags_453_reset = reset;
  assign tags_454_clock = clock;
  assign tags_454_reset = reset;
  assign tags_455_clock = clock;
  assign tags_455_reset = reset;
  assign tags_456_clock = clock;
  assign tags_456_reset = reset;
  assign tags_457_clock = clock;
  assign tags_457_reset = reset;
  assign tags_458_clock = clock;
  assign tags_458_reset = reset;
  assign tags_459_clock = clock;
  assign tags_459_reset = reset;
  assign tags_460_clock = clock;
  assign tags_460_reset = reset;
  assign tags_461_clock = clock;
  assign tags_461_reset = reset;
  assign tags_462_clock = clock;
  assign tags_462_reset = reset;
  assign tags_463_clock = clock;
  assign tags_463_reset = reset;
  assign tags_464_clock = clock;
  assign tags_464_reset = reset;
  assign tags_465_clock = clock;
  assign tags_465_reset = reset;
  assign tags_466_clock = clock;
  assign tags_466_reset = reset;
  assign tags_467_clock = clock;
  assign tags_467_reset = reset;
  assign tags_468_clock = clock;
  assign tags_468_reset = reset;
  assign tags_469_clock = clock;
  assign tags_469_reset = reset;
  assign tags_470_clock = clock;
  assign tags_470_reset = reset;
  assign tags_471_clock = clock;
  assign tags_471_reset = reset;
  assign tags_472_clock = clock;
  assign tags_472_reset = reset;
  assign tags_473_clock = clock;
  assign tags_473_reset = reset;
  assign tags_474_clock = clock;
  assign tags_474_reset = reset;
  assign tags_475_clock = clock;
  assign tags_475_reset = reset;
  assign tags_476_clock = clock;
  assign tags_476_reset = reset;
  assign tags_477_clock = clock;
  assign tags_477_reset = reset;
  assign tags_478_clock = clock;
  assign tags_478_reset = reset;
  assign tags_479_clock = clock;
  assign tags_479_reset = reset;
  assign tags_480_clock = clock;
  assign tags_480_reset = reset;
  assign tags_481_clock = clock;
  assign tags_481_reset = reset;
  assign tags_482_clock = clock;
  assign tags_482_reset = reset;
  assign tags_483_clock = clock;
  assign tags_483_reset = reset;
  assign tags_484_clock = clock;
  assign tags_484_reset = reset;
  assign tags_485_clock = clock;
  assign tags_485_reset = reset;
  assign tags_486_clock = clock;
  assign tags_486_reset = reset;
  assign tags_487_clock = clock;
  assign tags_487_reset = reset;
  assign tags_488_clock = clock;
  assign tags_488_reset = reset;
  assign tags_489_clock = clock;
  assign tags_489_reset = reset;
  assign tags_490_clock = clock;
  assign tags_490_reset = reset;
  assign tags_491_clock = clock;
  assign tags_491_reset = reset;
  assign tags_492_clock = clock;
  assign tags_492_reset = reset;
  assign tags_493_clock = clock;
  assign tags_493_reset = reset;
  assign tags_494_clock = clock;
  assign tags_494_reset = reset;
  assign tags_495_clock = clock;
  assign tags_495_reset = reset;
  assign tags_496_clock = clock;
  assign tags_496_reset = reset;
  assign tags_497_clock = clock;
  assign tags_497_reset = reset;
  assign tags_498_clock = clock;
  assign tags_498_reset = reset;
  assign tags_499_clock = clock;
  assign tags_499_reset = reset;
  assign tags_500_clock = clock;
  assign tags_500_reset = reset;
  assign tags_501_clock = clock;
  assign tags_501_reset = reset;
  assign tags_502_clock = clock;
  assign tags_502_reset = reset;
  assign tags_503_clock = clock;
  assign tags_503_reset = reset;
  assign tags_504_clock = clock;
  assign tags_504_reset = reset;
  assign tags_505_clock = clock;
  assign tags_505_reset = reset;
  assign tags_506_clock = clock;
  assign tags_506_reset = reset;
  assign tags_507_clock = clock;
  assign tags_507_reset = reset;
  assign tags_508_clock = clock;
  assign tags_508_reset = reset;
  assign tags_509_clock = clock;
  assign tags_509_reset = reset;
  assign tags_510_clock = clock;
  assign tags_510_reset = reset;
  assign tags_511_clock = clock;
  assign tags_511_reset = reset;
  assign metadata_io_wdata_0 = md_0;
  assign metadata_io_wdata_1 = md_1;
  assign metadata_io_wdata_2 = md_2;
  assign metadata_io_wdata_3 = md_3;
  assign metadata_io_wdata_4 = md_4;
  assign metadata_io_wdata_5 = md_5;
  assign metadata_io_wdata_6 = md_6;
  assign metadata_io_wdata_7 = md_7;
  assign metadata_io_wdata_8 = md_8;
  assign metadata_io_wdata_9 = md_9;
  assign metadata_io_wdata_10 = md_10;
  assign metadata_io_wdata_11 = md_11;
  assign metadata_io_wdata_12 = md_12;
  assign metadata_io_wdata_13 = md_13;
  assign metadata_io_wdata_14 = md_14;
  assign metadata_io_wdata_15 = md_15;
  assign metadata_clock = clock;
  assign woffset = _T_19089;
  assign md_0 = _GEN_2;
  assign md_1 = _GEN_3;
  assign md_2 = _GEN_4;
  assign md_3 = _GEN_5;
  assign md_4 = _GEN_6;
  assign md_5 = _GEN_7;
  assign md_6 = _GEN_8;
  assign md_7 = _GEN_9;
  assign md_8 = _GEN_10;
  assign md_9 = _GEN_11;
  assign md_10 = _GEN_12;
  assign md_11 = _GEN_13;
  assign md_12 = _GEN_14;
  assign md_13 = _GEN_15;
  assign md_14 = _GEN_16;
  assign md_15 = _GEN_17;
  assign _GEN_0 = {{3'd0}, _T_19127};
endmodule
module FIFOCounter(
  input   clock,
  input   reset,
  input   io_enqVld,
  output  io_full,
  output  io_almostFull
);
  wire  sizeUDC_clock;
  wire  sizeUDC_reset;
  wire [9:0] sizeUDC_io_strideInc;
  wire [9:0] sizeUDC_io_strideDec;
  wire  sizeUDC_io_dec;
  wire [9:0] sizeUDC_io_out;
  wire [9:0] sizeUDC_io_nextInc;
  wire [9:0] sizeUDC_io_nextDec;
  wire [10:0] _T_23;
  wire [10:0] _T_24;
  wire [9:0] remainingSlots;
  wire [10:0] _T_26;
  wire [10:0] _T_27;
  wire [9:0] nextRemainingSlots;
  wire  full;
  wire  almostFull;
  UpDownCtr sizeUDC (
    .clock(sizeUDC_clock),
    .reset(sizeUDC_reset),
    .io_strideInc(sizeUDC_io_strideInc),
    .io_strideDec(sizeUDC_io_strideDec),
    .io_dec(sizeUDC_io_dec),
    .io_out(sizeUDC_io_out),
    .io_nextInc(sizeUDC_io_nextInc),
    .io_nextDec(sizeUDC_io_nextDec)
  );
  assign _T_23 = 10'h200 - sizeUDC_io_out;
  assign _T_24 = $unsigned(_T_23);
  assign remainingSlots = _T_24[9:0];
  assign _T_26 = 10'h200 - sizeUDC_io_nextInc;
  assign _T_27 = $unsigned(_T_26);
  assign nextRemainingSlots = _T_27[9:0];
  assign full = remainingSlots < 10'h1;
  assign almostFull = nextRemainingSlots < 10'h1;
  assign io_full = full;
  assign io_almostFull = almostFull;
  assign sizeUDC_io_strideInc = 10'h1;
  assign sizeUDC_io_strideDec = 10'h1;
  assign sizeUDC_io_dec = 1'h0;
  assign sizeUDC_clock = clock;
  assign sizeUDC_reset = reset;
endmodule
module MuxNType_17(
  input   io_ins_0,
  output  io_out
);
  assign io_out = io_ins_0;
endmodule
module RetimeWrapper_1113(
  input         clock,
  input         reset,
  input  [39:0] io_in,
  output [39:0] io_out
);
  wire [39:0] sr_out;
  wire [39:0] sr_in;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_1114(
  input         clock,
  input         reset,
  input  [39:0] io_in,
  output [39:0] io_out,
  input         io_enable
);
  wire [39:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [39:0] RetimeWrapper_io_in;
  wire [39:0] RetimeWrapper_io_out;
  wire [39:0] _T_9;
  wire [39:0] _GEN_0;
  wire [39:0] _GEN_1;
  RetimeWrapper_1113 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? 40'h0 : _T_9;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_9;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_9 = RetimeWrapper_io_out;
endmodule
module Counter_19(
  input         clock,
  input         reset,
  input  [39:0] io_max,
  output [39:0] io_out,
  input         io_enable,
  input         io_saturate,
  output        io_done
);
  wire  reg$_clock;
  wire  reg$_reset;
  wire [39:0] reg$_io_in;
  wire [39:0] reg$_io_out;
  wire  reg$_io_enable;
  wire [40:0] count;
  wire [41:0] _T_12;
  wire [40:0] newval;
  wire [40:0] _GEN_1;
  wire  isMax;
  wire [40:0] _T_13;
  wire [40:0] next;
  wire  _T_14;
  FF_1114 reg$ (
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out};
  assign _T_12 = count + 41'h1;
  assign newval = _T_12[40:0];
  assign _GEN_1 = {{1'd0}, io_max};
  assign isMax = newval >= _GEN_1;
  assign _T_13 = io_saturate ? count : 41'h0;
  assign next = isMax ? _T_13 : newval;
  assign _T_14 = io_enable & isMax;
  assign io_out = count[39:0];
  assign io_done = _T_14;
  assign reg$_io_in = next[39:0];
  assign reg$_io_enable = io_enable;
  assign reg$_clock = clock;
  assign reg$_reset = reset;
endmodule
module RetimeWrapper_1159(
  input         clock,
  input         reset,
  input  [63:0] io_in,
  output [63:0] io_out
);
  wire [63:0] sr_out;
  wire [63:0] sr_in;
  wire  sr_reset;
  wire  sr_clock;
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr (
    .out(sr_out),
    .in(sr_in),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out;
  assign sr_in = io_in;
  assign sr_reset = reset;
  assign sr_clock = clock;
endmodule
module FF_1160(
  input         clock,
  input         reset,
  input  [63:0] io_in,
  input  [63:0] io_init,
  output [63:0] io_out,
  input         io_enable
);
  wire [63:0] d;
  wire  RetimeWrapper_clock;
  wire  RetimeWrapper_reset;
  wire [63:0] RetimeWrapper_io_in;
  wire [63:0] RetimeWrapper_io_out;
  wire [63:0] _T_9;
  wire [63:0] _GEN_0;
  wire [63:0] _GEN_1;
  RetimeWrapper_1159 RetimeWrapper (
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _GEN_0 = reset ? io_init : _T_9;
  assign _GEN_1 = io_enable ? io_in : _GEN_0;
  assign io_out = _T_9;
  assign d = _GEN_1;
  assign RetimeWrapper_io_in = d;
  assign RetimeWrapper_clock = clock;
  assign RetimeWrapper_reset = reset;
  assign _T_9 = RetimeWrapper_io_out;
endmodule
module MAGCore(
  input         clock,
  input         reset,
  input         io_enable,
  output [31:0] io_debugSignals_0,
  output [31:0] io_debugSignals_1,
  output [31:0] io_debugSignals_2,
  output [31:0] io_debugSignals_3,
  output [31:0] io_debugSignals_4,
  output [31:0] io_debugSignals_5,
  output [31:0] io_debugSignals_6,
  output [31:0] io_debugSignals_7,
  output [31:0] io_debugSignals_8,
  output [31:0] io_debugSignals_9,
  output [31:0] io_debugSignals_10,
  output [31:0] io_debugSignals_11,
  output [31:0] io_debugSignals_12,
  output [31:0] io_debugSignals_13,
  output [31:0] io_debugSignals_14,
  output [31:0] io_debugSignals_15,
  output [31:0] io_debugSignals_16,
  output [31:0] io_debugSignals_17,
  output [31:0] io_debugSignals_18,
  output [31:0] io_debugSignals_19,
  output [31:0] io_debugSignals_20,
  output [31:0] io_debugSignals_21,
  output [31:0] io_debugSignals_22,
  output [31:0] io_debugSignals_23,
  output [31:0] io_debugSignals_24,
  output [31:0] io_debugSignals_25,
  output [31:0] io_debugSignals_26,
  output [31:0] io_debugSignals_27,
  output [31:0] io_debugSignals_28,
  output [31:0] io_debugSignals_29,
  output [31:0] io_debugSignals_30,
  output [31:0] io_debugSignals_31,
  output [31:0] io_debugSignals_32,
  output [31:0] io_debugSignals_33,
  output [31:0] io_debugSignals_34,
  output [31:0] io_debugSignals_35,
  output [31:0] io_debugSignals_36,
  output [31:0] io_debugSignals_37,
  output [31:0] io_debugSignals_38,
  output [31:0] io_debugSignals_39,
  output [31:0] io_debugSignals_40,
  output [31:0] io_debugSignals_41,
  output [31:0] io_debugSignals_42,
  output [31:0] io_debugSignals_43,
  output [31:0] io_debugSignals_44,
  output [31:0] io_debugSignals_45,
  output [31:0] io_debugSignals_46,
  output [31:0] io_debugSignals_47,
  output [31:0] io_debugSignals_48,
  output [31:0] io_debugSignals_49,
  output [31:0] io_debugSignals_50,
  output [31:0] io_debugSignals_51,
  output [31:0] io_debugSignals_52,
  output [31:0] io_debugSignals_53,
  output [31:0] io_debugSignals_54,
  output [31:0] io_debugSignals_55,
  output [31:0] io_debugSignals_56,
  output [31:0] io_debugSignals_57,
  output [31:0] io_debugSignals_58,
  output        io_dram_rresp_ready
);
  wire  commandFifo_clock;
  wire  commandFifo_reset;
  wire [81:0] commandFifo_io_deq_0;
  wire  commandFifo_io_deqVld;
  wire  commandFifo_io_empty;
  wire  commandFifo_io_tag;
  wire [63:0] headCommand_addr;
  wire  headCommand_isWr;
  wire  headCommand_isSparse;
  wire [15:0] headCommand_size;
  wire [63:0] _T_484_addr;
  wire  _T_484_isWr;
  wire  _T_484_isSparse;
  wire [15:0] _T_484_size;
  wire [63:0] _T_485;
  wire  _T_486;
  wire  _T_487;
  wire [15:0] _T_488;
  wire  _T_495;
  wire  isSparse;
  wire [9:0] _T_497;
  wire [5:0] _T_498;
  wire  _T_500;
  wire [9:0] _GEN_0;
  wire [10:0] _T_501;
  wire [9:0] sizeInBursts;
  wire  wdataFifo_clock;
  wire  wdataFifo_reset;
  wire  wdataFifo_io_empty;
  wire  wdataFifo_io_forceTag_valid;
  wire  wdataFifo_io_forceTag_bits;
  wire  wrPhase_clock;
  wire  wrPhase_reset;
  wire  wrPhase_io_input_set;
  wire  wrPhase_io_input_reset;
  wire  wrPhase_io_input_asyn_reset;
  wire  wrPhase_io_output_data;
  wire  burstVld;
  wire  _T_506;
  wire  writeCmd;
  wire  _T_507;
  wire  wdataValid;
  wire [1:0] _T_509;
  wire [1:0] _T_510;
  wire  _T_511;
  wire  _T_513;
  wire  sparseWriteEnable;
  wire  _T_515;
  wire  _T_517;
  wire  issuedFF_clock;
  wire  issuedFF_reset;
  wire  issuedFF_io_in;
  wire  issuedFF_io_out;
  wire  issuedFF_io_enable;
  wire  burstCounter_clock;
  wire  burstCounter_reset;
  wire [31:0] burstCounter_io_max;
  wire [31:0] burstCounter_io_out;
  wire  burstCounter_io_enable;
  wire  burstCounter_io_done;
  wire [9:0] _T_525;
  wire  dramReadySeen;
  wire  dramReadyFF_clock;
  wire  dramReadyFF_reset;
  wire  dramReadyFF_io_in;
  wire  dramReadyFF_io_out;
  wire  dramReadyFF_io_enable;
  wire  _T_536;
  wire  _T_537;
  wire  _T_540;
  wire  _T_544;
  wire  _T_545;
  wire  _T_546;
  wire  _T_548;
  wire  _T_549;
  wire  burstTagCounter_clock;
  wire  burstTagCounter_reset;
  wire [10:0] burstTagCounter_io_out;
  wire [3:0] elementID;
  wire  wdataSelectCounter_clock;
  wire  wdataSelectCounter_reset;
  wire  wdataSelectCounter_io_reset;
  wire  _T_567;
  wire  ccache_clock;
  wire  ccache_reset;
  wire [7:0] ccache_io_rmetaData_0;
  wire [7:0] ccache_io_rmetaData_1;
  wire [7:0] ccache_io_rmetaData_2;
  wire [7:0] ccache_io_rmetaData_3;
  wire [7:0] ccache_io_rmetaData_4;
  wire [7:0] ccache_io_rmetaData_5;
  wire [7:0] ccache_io_rmetaData_6;
  wire [7:0] ccache_io_rmetaData_7;
  wire [7:0] ccache_io_rmetaData_8;
  wire [7:0] ccache_io_rmetaData_9;
  wire [7:0] ccache_io_rmetaData_10;
  wire [7:0] ccache_io_rmetaData_11;
  wire [7:0] ccache_io_rmetaData_12;
  wire [7:0] ccache_io_rmetaData_13;
  wire [7:0] ccache_io_rmetaData_14;
  wire [7:0] ccache_io_rmetaData_15;
  wire [31:0] ccache_io_waddr;
  wire [3:0] ccache_io_position;
  wire  sgValidDepulser_clock;
  wire  sgValidDepulser_reset;
  wire  sgValidDepulser_io_in;
  wire  sgValidDepulser_io_rst;
  wire  sgValidDepulser_io_out;
  wire  _T_580;
  wire  validMask_0;
  wire  validMask_1;
  wire  validMask_2;
  wire  validMask_3;
  wire  validMask_4;
  wire  validMask_5;
  wire  validMask_6;
  wire  validMask_7;
  wire  validMask_8;
  wire  validMask_9;
  wire  validMask_10;
  wire  validMask_11;
  wire  validMask_12;
  wire  validMask_13;
  wire  validMask_14;
  wire  validMask_15;
  wire  gatherBuffer_0_clock;
  wire  gatherBuffer_0_reset;
  wire [31:0] gatherBuffer_0_io_in;
  wire [31:0] gatherBuffer_0_io_init;
  wire [31:0] gatherBuffer_0_io_out;
  wire  gatherBuffer_0_io_enable;
  wire  gatherBuffer_1_clock;
  wire  gatherBuffer_1_reset;
  wire [31:0] gatherBuffer_1_io_in;
  wire [31:0] gatherBuffer_1_io_init;
  wire [31:0] gatherBuffer_1_io_out;
  wire  gatherBuffer_1_io_enable;
  wire  gatherBuffer_2_clock;
  wire  gatherBuffer_2_reset;
  wire [31:0] gatherBuffer_2_io_in;
  wire [31:0] gatherBuffer_2_io_init;
  wire [31:0] gatherBuffer_2_io_out;
  wire  gatherBuffer_2_io_enable;
  wire  gatherBuffer_3_clock;
  wire  gatherBuffer_3_reset;
  wire [31:0] gatherBuffer_3_io_in;
  wire [31:0] gatherBuffer_3_io_init;
  wire [31:0] gatherBuffer_3_io_out;
  wire  gatherBuffer_3_io_enable;
  wire  gatherBuffer_4_clock;
  wire  gatherBuffer_4_reset;
  wire [31:0] gatherBuffer_4_io_in;
  wire [31:0] gatherBuffer_4_io_init;
  wire [31:0] gatherBuffer_4_io_out;
  wire  gatherBuffer_4_io_enable;
  wire  gatherBuffer_5_clock;
  wire  gatherBuffer_5_reset;
  wire [31:0] gatherBuffer_5_io_in;
  wire [31:0] gatherBuffer_5_io_init;
  wire [31:0] gatherBuffer_5_io_out;
  wire  gatherBuffer_5_io_enable;
  wire  gatherBuffer_6_clock;
  wire  gatherBuffer_6_reset;
  wire [31:0] gatherBuffer_6_io_in;
  wire [31:0] gatherBuffer_6_io_init;
  wire [31:0] gatherBuffer_6_io_out;
  wire  gatherBuffer_6_io_enable;
  wire  gatherBuffer_7_clock;
  wire  gatherBuffer_7_reset;
  wire [31:0] gatherBuffer_7_io_in;
  wire [31:0] gatherBuffer_7_io_init;
  wire [31:0] gatherBuffer_7_io_out;
  wire  gatherBuffer_7_io_enable;
  wire  gatherBuffer_8_clock;
  wire  gatherBuffer_8_reset;
  wire [31:0] gatherBuffer_8_io_in;
  wire [31:0] gatherBuffer_8_io_init;
  wire [31:0] gatherBuffer_8_io_out;
  wire  gatherBuffer_8_io_enable;
  wire  gatherBuffer_9_clock;
  wire  gatherBuffer_9_reset;
  wire [31:0] gatherBuffer_9_io_in;
  wire [31:0] gatherBuffer_9_io_init;
  wire [31:0] gatherBuffer_9_io_out;
  wire  gatherBuffer_9_io_enable;
  wire  gatherBuffer_10_clock;
  wire  gatherBuffer_10_reset;
  wire [31:0] gatherBuffer_10_io_in;
  wire [31:0] gatherBuffer_10_io_init;
  wire [31:0] gatherBuffer_10_io_out;
  wire  gatherBuffer_10_io_enable;
  wire  gatherBuffer_11_clock;
  wire  gatherBuffer_11_reset;
  wire [31:0] gatherBuffer_11_io_in;
  wire [31:0] gatherBuffer_11_io_init;
  wire [31:0] gatherBuffer_11_io_out;
  wire  gatherBuffer_11_io_enable;
  wire  gatherBuffer_12_clock;
  wire  gatherBuffer_12_reset;
  wire [31:0] gatherBuffer_12_io_in;
  wire [31:0] gatherBuffer_12_io_init;
  wire [31:0] gatherBuffer_12_io_out;
  wire  gatherBuffer_12_io_enable;
  wire  gatherBuffer_13_clock;
  wire  gatherBuffer_13_reset;
  wire [31:0] gatherBuffer_13_io_in;
  wire [31:0] gatherBuffer_13_io_init;
  wire [31:0] gatherBuffer_13_io_out;
  wire  gatherBuffer_13_io_enable;
  wire  gatherBuffer_14_clock;
  wire  gatherBuffer_14_reset;
  wire [31:0] gatherBuffer_14_io_in;
  wire [31:0] gatherBuffer_14_io_init;
  wire [31:0] gatherBuffer_14_io_out;
  wire  gatherBuffer_14_io_enable;
  wire  gatherBuffer_15_clock;
  wire  gatherBuffer_15_reset;
  wire [31:0] gatherBuffer_15_io_in;
  wire [31:0] gatherBuffer_15_io_init;
  wire [31:0] gatherBuffer_15_io_out;
  wire  gatherBuffer_15_io_enable;
  wire  completionMask_0_clock;
  wire  completionMask_0_reset;
  wire  completionMask_0_io_in;
  wire  completionMask_0_io_out;
  wire  completionMask_0_io_enable;
  wire  completionMask_1_clock;
  wire  completionMask_1_reset;
  wire  completionMask_1_io_in;
  wire  completionMask_1_io_out;
  wire  completionMask_1_io_enable;
  wire  completionMask_2_clock;
  wire  completionMask_2_reset;
  wire  completionMask_2_io_in;
  wire  completionMask_2_io_out;
  wire  completionMask_2_io_enable;
  wire  completionMask_3_clock;
  wire  completionMask_3_reset;
  wire  completionMask_3_io_in;
  wire  completionMask_3_io_out;
  wire  completionMask_3_io_enable;
  wire  completionMask_4_clock;
  wire  completionMask_4_reset;
  wire  completionMask_4_io_in;
  wire  completionMask_4_io_out;
  wire  completionMask_4_io_enable;
  wire  completionMask_5_clock;
  wire  completionMask_5_reset;
  wire  completionMask_5_io_in;
  wire  completionMask_5_io_out;
  wire  completionMask_5_io_enable;
  wire  completionMask_6_clock;
  wire  completionMask_6_reset;
  wire  completionMask_6_io_in;
  wire  completionMask_6_io_out;
  wire  completionMask_6_io_enable;
  wire  completionMask_7_clock;
  wire  completionMask_7_reset;
  wire  completionMask_7_io_in;
  wire  completionMask_7_io_out;
  wire  completionMask_7_io_enable;
  wire  completionMask_8_clock;
  wire  completionMask_8_reset;
  wire  completionMask_8_io_in;
  wire  completionMask_8_io_out;
  wire  completionMask_8_io_enable;
  wire  completionMask_9_clock;
  wire  completionMask_9_reset;
  wire  completionMask_9_io_in;
  wire  completionMask_9_io_out;
  wire  completionMask_9_io_enable;
  wire  completionMask_10_clock;
  wire  completionMask_10_reset;
  wire  completionMask_10_io_in;
  wire  completionMask_10_io_out;
  wire  completionMask_10_io_enable;
  wire  completionMask_11_clock;
  wire  completionMask_11_reset;
  wire  completionMask_11_io_in;
  wire  completionMask_11_io_out;
  wire  completionMask_11_io_enable;
  wire  completionMask_12_clock;
  wire  completionMask_12_reset;
  wire  completionMask_12_io_in;
  wire  completionMask_12_io_out;
  wire  completionMask_12_io_enable;
  wire  completionMask_13_clock;
  wire  completionMask_13_reset;
  wire  completionMask_13_io_in;
  wire  completionMask_13_io_out;
  wire  completionMask_13_io_enable;
  wire  completionMask_14_clock;
  wire  completionMask_14_reset;
  wire  completionMask_14_io_in;
  wire  completionMask_14_io_out;
  wire  completionMask_14_io_enable;
  wire  completionMask_15_clock;
  wire  completionMask_15_reset;
  wire  completionMask_15_io_in;
  wire  completionMask_15_io_out;
  wire  completionMask_15_io_enable;
  wire [10:0] _T_845;
  wire [10:0] _T_846;
  wire [9:0] _T_847;
  wire [31:0] _GEN_1;
  wire  _T_848;
  wire  wlast;
  wire  wasSparseWren_clock;
  wire  wasSparseWren_reset;
  wire  wasSparseWren_io_input_set;
  wire  wasSparseWren_io_input_reset;
  wire  wasSparseWren_io_input_asyn_reset;
  wire  wasSparseWren_io_output_data;
  wire  _T_849;
  wire  _T_852;
  wire  _T_853;
  reg  _T_856;
  reg [31:0] _RAND_0;
  wire  rdataFifos_0_clock;
  wire  rdataFifos_0_reset;
  wire  rdataFifos_0_io_enqVld;
  wire  rdataFifos_0_io_full;
  wire  rdataFifos_0_io_empty;
  wire  rdataFifos_0_io_almostFull;
  wire  _T_869;
  wire  _T_870;
  wire  wrespFifos_0_clock;
  wire  wrespFifos_0_reset;
  wire  wrespFifos_0_io_enqVld;
  wire  wrespFifos_0_io_full;
  wire  wrespFifos_0_io_almostFull;
  wire  MuxNType_1_io_ins_0;
  wire  MuxNType_1_io_out;
  wire  _T_886_0;
  wire  MuxNType_2_io_ins_0;
  wire  MuxNType_2_io_out;
  wire  _T_890;
  wire  _T_891;
  wire  _T_894_0;
  wire  Counter_clock;
  wire  Counter_reset;
  wire [39:0] Counter_io_max;
  wire [39:0] Counter_io_out;
  wire  Counter_io_enable;
  wire  Counter_io_saturate;
  wire  Counter_io_done;
  wire  Counter_1_clock;
  wire  Counter_1_reset;
  wire [31:0] Counter_1_io_max;
  wire [31:0] Counter_1_io_out;
  wire  Counter_1_io_enable;
  wire  Counter_1_io_done;
  wire  FF_clock;
  wire  FF_reset;
  wire [31:0] FF_io_in;
  wire [31:0] FF_io_init;
  wire [31:0] FF_io_out;
  wire  FF_io_enable;
  wire  FF_1_clock;
  wire  FF_1_reset;
  wire [31:0] FF_1_io_in;
  wire [31:0] FF_1_io_init;
  wire [31:0] FF_1_io_out;
  wire  FF_1_io_enable;
  wire  FF_2_clock;
  wire  FF_2_reset;
  wire [31:0] FF_2_io_in;
  wire [31:0] FF_2_io_init;
  wire [31:0] FF_2_io_out;
  wire  FF_2_io_enable;
  wire  FF_3_clock;
  wire  FF_3_reset;
  wire [31:0] FF_3_io_in;
  wire [31:0] FF_3_io_init;
  wire [31:0] FF_3_io_out;
  wire  FF_3_io_enable;
  wire  FF_4_clock;
  wire  FF_4_reset;
  wire [31:0] FF_4_io_in;
  wire [31:0] FF_4_io_init;
  wire [31:0] FF_4_io_out;
  wire  FF_4_io_enable;
  wire  FF_5_clock;
  wire  FF_5_reset;
  wire [31:0] FF_5_io_in;
  wire [31:0] FF_5_io_init;
  wire [31:0] FF_5_io_out;
  wire  FF_5_io_enable;
  wire  FF_6_clock;
  wire  FF_6_reset;
  wire [31:0] FF_6_io_in;
  wire [31:0] FF_6_io_init;
  wire [31:0] FF_6_io_out;
  wire  FF_6_io_enable;
  wire  FF_7_clock;
  wire  FF_7_reset;
  wire [31:0] FF_7_io_in;
  wire [31:0] FF_7_io_init;
  wire [31:0] FF_7_io_out;
  wire  FF_7_io_enable;
  wire  FF_8_clock;
  wire  FF_8_reset;
  wire [31:0] FF_8_io_in;
  wire [31:0] FF_8_io_init;
  wire [31:0] FF_8_io_out;
  wire  FF_8_io_enable;
  wire  FF_9_clock;
  wire  FF_9_reset;
  wire [31:0] FF_9_io_in;
  wire [31:0] FF_9_io_init;
  wire [31:0] FF_9_io_out;
  wire  FF_9_io_enable;
  wire  FF_10_clock;
  wire  FF_10_reset;
  wire [31:0] FF_10_io_in;
  wire [31:0] FF_10_io_init;
  wire [31:0] FF_10_io_out;
  wire  FF_10_io_enable;
  wire  FF_11_clock;
  wire  FF_11_reset;
  wire [31:0] FF_11_io_in;
  wire [31:0] FF_11_io_init;
  wire [31:0] FF_11_io_out;
  wire  FF_11_io_enable;
  wire  FF_12_clock;
  wire  FF_12_reset;
  wire [31:0] FF_12_io_in;
  wire [31:0] FF_12_io_init;
  wire [31:0] FF_12_io_out;
  wire  FF_12_io_enable;
  wire  FF_13_clock;
  wire  FF_13_reset;
  wire [31:0] FF_13_io_in;
  wire [31:0] FF_13_io_init;
  wire [31:0] FF_13_io_out;
  wire  FF_13_io_enable;
  wire  FF_14_clock;
  wire  FF_14_reset;
  wire [31:0] FF_14_io_in;
  wire [31:0] FF_14_io_init;
  wire [31:0] FF_14_io_out;
  wire  FF_14_io_enable;
  wire  FF_15_clock;
  wire  FF_15_reset;
  wire [31:0] FF_15_io_in;
  wire [31:0] FF_15_io_init;
  wire [31:0] FF_15_io_out;
  wire  FF_15_io_enable;
  wire  FF_16_clock;
  wire  FF_16_reset;
  wire [31:0] FF_16_io_in;
  wire [31:0] FF_16_io_init;
  wire [31:0] FF_16_io_out;
  wire  FF_16_io_enable;
  wire  FF_17_clock;
  wire  FF_17_reset;
  wire [31:0] FF_17_io_in;
  wire [31:0] FF_17_io_init;
  wire [31:0] FF_17_io_out;
  wire  FF_17_io_enable;
  wire  FF_18_clock;
  wire  FF_18_reset;
  wire [31:0] FF_18_io_in;
  wire [31:0] FF_18_io_init;
  wire [31:0] FF_18_io_out;
  wire  FF_18_io_enable;
  wire  FF_19_clock;
  wire  FF_19_reset;
  wire [31:0] FF_19_io_in;
  wire [31:0] FF_19_io_init;
  wire [31:0] FF_19_io_out;
  wire  FF_19_io_enable;
  wire  FF_20_clock;
  wire  FF_20_reset;
  wire [31:0] FF_20_io_in;
  wire [31:0] FF_20_io_init;
  wire [31:0] FF_20_io_out;
  wire  FF_20_io_enable;
  wire  FF_21_clock;
  wire  FF_21_reset;
  wire [31:0] FF_21_io_in;
  wire [31:0] FF_21_io_init;
  wire [31:0] FF_21_io_out;
  wire  FF_21_io_enable;
  wire  FF_22_clock;
  wire  FF_22_reset;
  wire [31:0] FF_22_io_in;
  wire [31:0] FF_22_io_init;
  wire [31:0] FF_22_io_out;
  wire  FF_22_io_enable;
  wire  FF_23_clock;
  wire  FF_23_reset;
  wire [31:0] FF_23_io_in;
  wire [31:0] FF_23_io_init;
  wire [31:0] FF_23_io_out;
  wire  FF_23_io_enable;
  wire  FF_24_clock;
  wire  FF_24_reset;
  wire [31:0] FF_24_io_in;
  wire [31:0] FF_24_io_init;
  wire [31:0] FF_24_io_out;
  wire  FF_24_io_enable;
  wire  FF_25_clock;
  wire  FF_25_reset;
  wire [31:0] FF_25_io_in;
  wire [31:0] FF_25_io_init;
  wire [31:0] FF_25_io_out;
  wire  FF_25_io_enable;
  wire  FF_26_clock;
  wire  FF_26_reset;
  wire [31:0] FF_26_io_in;
  wire [31:0] FF_26_io_init;
  wire [31:0] FF_26_io_out;
  wire  FF_26_io_enable;
  wire  FF_27_clock;
  wire  FF_27_reset;
  wire [31:0] FF_27_io_in;
  wire [31:0] FF_27_io_init;
  wire [31:0] FF_27_io_out;
  wire  FF_27_io_enable;
  wire  FF_28_clock;
  wire  FF_28_reset;
  wire [31:0] FF_28_io_in;
  wire [31:0] FF_28_io_init;
  wire [31:0] FF_28_io_out;
  wire  FF_28_io_enable;
  wire  FF_29_clock;
  wire  FF_29_reset;
  wire [31:0] FF_29_io_in;
  wire [31:0] FF_29_io_init;
  wire [31:0] FF_29_io_out;
  wire  FF_29_io_enable;
  wire  FF_30_clock;
  wire  FF_30_reset;
  wire [31:0] FF_30_io_in;
  wire [31:0] FF_30_io_init;
  wire [31:0] FF_30_io_out;
  wire  FF_30_io_enable;
  wire  FF_31_clock;
  wire  FF_31_reset;
  wire [31:0] FF_31_io_in;
  wire [31:0] FF_31_io_init;
  wire [31:0] FF_31_io_out;
  wire  FF_31_io_enable;
  wire  Counter_2_clock;
  wire  Counter_2_reset;
  wire [31:0] Counter_2_io_max;
  wire [31:0] Counter_2_io_out;
  wire  Counter_2_io_enable;
  wire  Counter_2_io_done;
  wire  Counter_3_clock;
  wire  Counter_3_reset;
  wire [31:0] Counter_3_io_max;
  wire [31:0] Counter_3_io_out;
  wire  Counter_3_io_enable;
  wire  Counter_3_io_done;
  wire  Counter_4_clock;
  wire  Counter_4_reset;
  wire [31:0] Counter_4_io_max;
  wire [31:0] Counter_4_io_out;
  wire  Counter_4_io_enable;
  wire  Counter_4_io_done;
  wire  Counter_5_clock;
  wire  Counter_5_reset;
  wire [31:0] Counter_5_io_max;
  wire [31:0] Counter_5_io_out;
  wire  Counter_5_io_enable;
  wire  Counter_5_io_done;
  wire  Counter_6_clock;
  wire  Counter_6_reset;
  wire [31:0] Counter_6_io_max;
  wire [31:0] Counter_6_io_out;
  wire  Counter_6_io_enable;
  wire  Counter_6_io_done;
  wire  Counter_7_clock;
  wire  Counter_7_reset;
  wire [31:0] Counter_7_io_max;
  wire [31:0] Counter_7_io_out;
  wire  Counter_7_io_enable;
  wire  Counter_7_io_done;
  wire  Counter_8_clock;
  wire  Counter_8_reset;
  wire [31:0] Counter_8_io_max;
  wire [31:0] Counter_8_io_out;
  wire  Counter_8_io_enable;
  wire  Counter_8_io_done;
  wire  Counter_9_clock;
  wire  Counter_9_reset;
  wire [31:0] Counter_9_io_max;
  wire [31:0] Counter_9_io_out;
  wire  Counter_9_io_enable;
  wire  Counter_9_io_done;
  wire  Counter_10_clock;
  wire  Counter_10_reset;
  wire [31:0] Counter_10_io_max;
  wire [31:0] Counter_10_io_out;
  wire  Counter_10_io_enable;
  wire  Counter_10_io_done;
  wire  Counter_11_clock;
  wire  Counter_11_reset;
  wire [31:0] Counter_11_io_max;
  wire [31:0] Counter_11_io_out;
  wire  Counter_11_io_enable;
  wire  Counter_11_io_done;
  wire  Counter_12_clock;
  wire  Counter_12_reset;
  wire [31:0] Counter_12_io_max;
  wire [31:0] Counter_12_io_out;
  wire  Counter_12_io_enable;
  wire  Counter_12_io_done;
  wire  Counter_13_clock;
  wire  Counter_13_reset;
  wire [31:0] Counter_13_io_max;
  wire [31:0] Counter_13_io_out;
  wire  Counter_13_io_enable;
  wire  Counter_13_io_done;
  wire  FF_32_clock;
  wire  FF_32_reset;
  wire [63:0] FF_32_io_in;
  wire [63:0] FF_32_io_init;
  wire [63:0] FF_32_io_out;
  wire  FF_32_io_enable;
  wire  FF_33_clock;
  wire  FF_33_reset;
  wire [63:0] FF_33_io_in;
  wire [63:0] FF_33_io_init;
  wire [63:0] FF_33_io_out;
  wire  FF_33_io_enable;
  wire  Counter_14_clock;
  wire  Counter_14_reset;
  wire [31:0] Counter_14_io_max;
  wire [31:0] Counter_14_io_out;
  wire  Counter_14_io_enable;
  wire  Counter_14_io_done;
  wire  Counter_15_clock;
  wire  Counter_15_reset;
  wire [31:0] Counter_15_io_max;
  wire [31:0] Counter_15_io_out;
  wire  Counter_15_io_enable;
  wire  Counter_15_io_done;
  wire  _T_1241;
  wire  Counter_16_clock;
  wire  Counter_16_reset;
  wire [31:0] Counter_16_io_max;
  wire [31:0] Counter_16_io_out;
  wire  Counter_16_io_enable;
  wire  Counter_16_io_done;
  wire  _T_1249;
  wire  Counter_17_clock;
  wire  Counter_17_reset;
  wire [31:0] Counter_17_io_max;
  wire [31:0] Counter_17_io_out;
  wire  Counter_17_io_enable;
  wire  Counter_17_io_done;
  wire  _T_1257;
  wire  Counter_18_clock;
  wire  Counter_18_reset;
  wire [31:0] Counter_18_io_max;
  wire [31:0] Counter_18_io_out;
  wire  Counter_18_io_enable;
  wire  Counter_18_io_done;
  wire  Counter_19_clock;
  wire  Counter_19_reset;
  wire [31:0] Counter_19_io_max;
  wire [31:0] Counter_19_io_out;
  wire  Counter_19_io_enable;
  wire  Counter_19_io_done;
  wire  Counter_20_clock;
  wire  Counter_20_reset;
  wire [31:0] Counter_20_io_max;
  wire [31:0] Counter_20_io_out;
  wire  Counter_20_io_enable;
  wire  Counter_20_io_done;
  wire  Counter_21_clock;
  wire  Counter_21_reset;
  wire [31:0] Counter_21_io_max;
  wire [31:0] Counter_21_io_out;
  wire  Counter_21_io_enable;
  wire  Counter_21_io_done;
  wire  Counter_22_clock;
  wire  Counter_22_reset;
  wire [31:0] Counter_22_io_max;
  wire [31:0] Counter_22_io_out;
  wire  Counter_22_io_enable;
  wire  Counter_22_io_done;
  wire  Counter_23_clock;
  wire  Counter_23_reset;
  wire [31:0] Counter_23_io_max;
  wire [31:0] Counter_23_io_out;
  wire  Counter_23_io_enable;
  wire  Counter_23_io_done;
  wire  Counter_24_clock;
  wire  Counter_24_reset;
  wire [31:0] Counter_24_io_max;
  wire [31:0] Counter_24_io_out;
  wire  Counter_24_io_enable;
  wire  Counter_24_io_done;
  wire  Counter_25_clock;
  wire  Counter_25_reset;
  wire [31:0] Counter_25_io_max;
  wire [31:0] Counter_25_io_out;
  wire  Counter_25_io_enable;
  wire  Counter_25_io_done;
  wire  Counter_26_clock;
  wire  Counter_26_reset;
  wire [31:0] Counter_26_io_max;
  wire [31:0] Counter_26_io_out;
  wire  Counter_26_io_enable;
  wire  Counter_26_io_done;
  FIFOArbiter commandFifo (
    .clock(commandFifo_clock),
    .reset(commandFifo_reset),
    .io_deq_0(commandFifo_io_deq_0),
    .io_deqVld(commandFifo_io_deqVld),
    .io_empty(commandFifo_io_empty),
    .io_tag(commandFifo_io_tag)
  );
  FIFOArbiterWidthConvert wdataFifo (
    .clock(wdataFifo_clock),
    .reset(wdataFifo_reset),
    .io_empty(wdataFifo_io_empty),
    .io_forceTag_valid(wdataFifo_io_forceTag_valid),
    .io_forceTag_bits(wdataFifo_io_forceTag_bits)
  );
  SRFF_sp wrPhase (
    .clock(wrPhase_clock),
    .reset(wrPhase_reset),
    .io_input_set(wrPhase_io_input_set),
    .io_input_reset(wrPhase_io_input_reset),
    .io_input_asyn_reset(wrPhase_io_input_asyn_reset),
    .io_output_data(wrPhase_io_output_data)
  );
  FF_9 issuedFF (
    .clock(issuedFF_clock),
    .reset(issuedFF_reset),
    .io_in(issuedFF_io_in),
    .io_out(issuedFF_io_out),
    .io_enable(issuedFF_io_enable)
  );
  Counter_12 burstCounter (
    .clock(burstCounter_clock),
    .reset(burstCounter_reset),
    .io_max(burstCounter_io_max),
    .io_out(burstCounter_io_out),
    .io_enable(burstCounter_io_enable),
    .io_done(burstCounter_io_done)
  );
  FF_9 dramReadyFF (
    .clock(dramReadyFF_clock),
    .reset(dramReadyFF_reset),
    .io_in(dramReadyFF_io_in),
    .io_out(dramReadyFF_io_out),
    .io_enable(dramReadyFF_io_enable)
  );
  Counter_13 burstTagCounter (
    .clock(burstTagCounter_clock),
    .reset(burstTagCounter_reset),
    .io_out(burstTagCounter_io_out)
  );
  Counter_14 wdataSelectCounter (
    .clock(wdataSelectCounter_clock),
    .reset(wdataSelectCounter_reset),
    .io_reset(wdataSelectCounter_io_reset)
  );
  CoalescingCache ccache (
    .clock(ccache_clock),
    .reset(ccache_reset),
    .io_rmetaData_0(ccache_io_rmetaData_0),
    .io_rmetaData_1(ccache_io_rmetaData_1),
    .io_rmetaData_2(ccache_io_rmetaData_2),
    .io_rmetaData_3(ccache_io_rmetaData_3),
    .io_rmetaData_4(ccache_io_rmetaData_4),
    .io_rmetaData_5(ccache_io_rmetaData_5),
    .io_rmetaData_6(ccache_io_rmetaData_6),
    .io_rmetaData_7(ccache_io_rmetaData_7),
    .io_rmetaData_8(ccache_io_rmetaData_8),
    .io_rmetaData_9(ccache_io_rmetaData_9),
    .io_rmetaData_10(ccache_io_rmetaData_10),
    .io_rmetaData_11(ccache_io_rmetaData_11),
    .io_rmetaData_12(ccache_io_rmetaData_12),
    .io_rmetaData_13(ccache_io_rmetaData_13),
    .io_rmetaData_14(ccache_io_rmetaData_14),
    .io_rmetaData_15(ccache_io_rmetaData_15),
    .io_waddr(ccache_io_waddr),
    .io_position(ccache_io_position)
  );
  Depulser sgValidDepulser (
    .clock(sgValidDepulser_clock),
    .reset(sgValidDepulser_reset),
    .io_in(sgValidDepulser_io_in),
    .io_rst(sgValidDepulser_io_rst),
    .io_out(sgValidDepulser_io_out)
  );
  FF_42 gatherBuffer_0 (
    .clock(gatherBuffer_0_clock),
    .reset(gatherBuffer_0_reset),
    .io_in(gatherBuffer_0_io_in),
    .io_init(gatherBuffer_0_io_init),
    .io_out(gatherBuffer_0_io_out),
    .io_enable(gatherBuffer_0_io_enable)
  );
  FF_42 gatherBuffer_1 (
    .clock(gatherBuffer_1_clock),
    .reset(gatherBuffer_1_reset),
    .io_in(gatherBuffer_1_io_in),
    .io_init(gatherBuffer_1_io_init),
    .io_out(gatherBuffer_1_io_out),
    .io_enable(gatherBuffer_1_io_enable)
  );
  FF_42 gatherBuffer_2 (
    .clock(gatherBuffer_2_clock),
    .reset(gatherBuffer_2_reset),
    .io_in(gatherBuffer_2_io_in),
    .io_init(gatherBuffer_2_io_init),
    .io_out(gatherBuffer_2_io_out),
    .io_enable(gatherBuffer_2_io_enable)
  );
  FF_42 gatherBuffer_3 (
    .clock(gatherBuffer_3_clock),
    .reset(gatherBuffer_3_reset),
    .io_in(gatherBuffer_3_io_in),
    .io_init(gatherBuffer_3_io_init),
    .io_out(gatherBuffer_3_io_out),
    .io_enable(gatherBuffer_3_io_enable)
  );
  FF_42 gatherBuffer_4 (
    .clock(gatherBuffer_4_clock),
    .reset(gatherBuffer_4_reset),
    .io_in(gatherBuffer_4_io_in),
    .io_init(gatherBuffer_4_io_init),
    .io_out(gatherBuffer_4_io_out),
    .io_enable(gatherBuffer_4_io_enable)
  );
  FF_42 gatherBuffer_5 (
    .clock(gatherBuffer_5_clock),
    .reset(gatherBuffer_5_reset),
    .io_in(gatherBuffer_5_io_in),
    .io_init(gatherBuffer_5_io_init),
    .io_out(gatherBuffer_5_io_out),
    .io_enable(gatherBuffer_5_io_enable)
  );
  FF_42 gatherBuffer_6 (
    .clock(gatherBuffer_6_clock),
    .reset(gatherBuffer_6_reset),
    .io_in(gatherBuffer_6_io_in),
    .io_init(gatherBuffer_6_io_init),
    .io_out(gatherBuffer_6_io_out),
    .io_enable(gatherBuffer_6_io_enable)
  );
  FF_42 gatherBuffer_7 (
    .clock(gatherBuffer_7_clock),
    .reset(gatherBuffer_7_reset),
    .io_in(gatherBuffer_7_io_in),
    .io_init(gatherBuffer_7_io_init),
    .io_out(gatherBuffer_7_io_out),
    .io_enable(gatherBuffer_7_io_enable)
  );
  FF_42 gatherBuffer_8 (
    .clock(gatherBuffer_8_clock),
    .reset(gatherBuffer_8_reset),
    .io_in(gatherBuffer_8_io_in),
    .io_init(gatherBuffer_8_io_init),
    .io_out(gatherBuffer_8_io_out),
    .io_enable(gatherBuffer_8_io_enable)
  );
  FF_42 gatherBuffer_9 (
    .clock(gatherBuffer_9_clock),
    .reset(gatherBuffer_9_reset),
    .io_in(gatherBuffer_9_io_in),
    .io_init(gatherBuffer_9_io_init),
    .io_out(gatherBuffer_9_io_out),
    .io_enable(gatherBuffer_9_io_enable)
  );
  FF_42 gatherBuffer_10 (
    .clock(gatherBuffer_10_clock),
    .reset(gatherBuffer_10_reset),
    .io_in(gatherBuffer_10_io_in),
    .io_init(gatherBuffer_10_io_init),
    .io_out(gatherBuffer_10_io_out),
    .io_enable(gatherBuffer_10_io_enable)
  );
  FF_42 gatherBuffer_11 (
    .clock(gatherBuffer_11_clock),
    .reset(gatherBuffer_11_reset),
    .io_in(gatherBuffer_11_io_in),
    .io_init(gatherBuffer_11_io_init),
    .io_out(gatherBuffer_11_io_out),
    .io_enable(gatherBuffer_11_io_enable)
  );
  FF_42 gatherBuffer_12 (
    .clock(gatherBuffer_12_clock),
    .reset(gatherBuffer_12_reset),
    .io_in(gatherBuffer_12_io_in),
    .io_init(gatherBuffer_12_io_init),
    .io_out(gatherBuffer_12_io_out),
    .io_enable(gatherBuffer_12_io_enable)
  );
  FF_42 gatherBuffer_13 (
    .clock(gatherBuffer_13_clock),
    .reset(gatherBuffer_13_reset),
    .io_in(gatherBuffer_13_io_in),
    .io_init(gatherBuffer_13_io_init),
    .io_out(gatherBuffer_13_io_out),
    .io_enable(gatherBuffer_13_io_enable)
  );
  FF_42 gatherBuffer_14 (
    .clock(gatherBuffer_14_clock),
    .reset(gatherBuffer_14_reset),
    .io_in(gatherBuffer_14_io_in),
    .io_init(gatherBuffer_14_io_init),
    .io_out(gatherBuffer_14_io_out),
    .io_enable(gatherBuffer_14_io_enable)
  );
  FF_42 gatherBuffer_15 (
    .clock(gatherBuffer_15_clock),
    .reset(gatherBuffer_15_reset),
    .io_in(gatherBuffer_15_io_in),
    .io_init(gatherBuffer_15_io_init),
    .io_out(gatherBuffer_15_io_out),
    .io_enable(gatherBuffer_15_io_enable)
  );
  FF_9 completionMask_0 (
    .clock(completionMask_0_clock),
    .reset(completionMask_0_reset),
    .io_in(completionMask_0_io_in),
    .io_out(completionMask_0_io_out),
    .io_enable(completionMask_0_io_enable)
  );
  FF_9 completionMask_1 (
    .clock(completionMask_1_clock),
    .reset(completionMask_1_reset),
    .io_in(completionMask_1_io_in),
    .io_out(completionMask_1_io_out),
    .io_enable(completionMask_1_io_enable)
  );
  FF_9 completionMask_2 (
    .clock(completionMask_2_clock),
    .reset(completionMask_2_reset),
    .io_in(completionMask_2_io_in),
    .io_out(completionMask_2_io_out),
    .io_enable(completionMask_2_io_enable)
  );
  FF_9 completionMask_3 (
    .clock(completionMask_3_clock),
    .reset(completionMask_3_reset),
    .io_in(completionMask_3_io_in),
    .io_out(completionMask_3_io_out),
    .io_enable(completionMask_3_io_enable)
  );
  FF_9 completionMask_4 (
    .clock(completionMask_4_clock),
    .reset(completionMask_4_reset),
    .io_in(completionMask_4_io_in),
    .io_out(completionMask_4_io_out),
    .io_enable(completionMask_4_io_enable)
  );
  FF_9 completionMask_5 (
    .clock(completionMask_5_clock),
    .reset(completionMask_5_reset),
    .io_in(completionMask_5_io_in),
    .io_out(completionMask_5_io_out),
    .io_enable(completionMask_5_io_enable)
  );
  FF_9 completionMask_6 (
    .clock(completionMask_6_clock),
    .reset(completionMask_6_reset),
    .io_in(completionMask_6_io_in),
    .io_out(completionMask_6_io_out),
    .io_enable(completionMask_6_io_enable)
  );
  FF_9 completionMask_7 (
    .clock(completionMask_7_clock),
    .reset(completionMask_7_reset),
    .io_in(completionMask_7_io_in),
    .io_out(completionMask_7_io_out),
    .io_enable(completionMask_7_io_enable)
  );
  FF_9 completionMask_8 (
    .clock(completionMask_8_clock),
    .reset(completionMask_8_reset),
    .io_in(completionMask_8_io_in),
    .io_out(completionMask_8_io_out),
    .io_enable(completionMask_8_io_enable)
  );
  FF_9 completionMask_9 (
    .clock(completionMask_9_clock),
    .reset(completionMask_9_reset),
    .io_in(completionMask_9_io_in),
    .io_out(completionMask_9_io_out),
    .io_enable(completionMask_9_io_enable)
  );
  FF_9 completionMask_10 (
    .clock(completionMask_10_clock),
    .reset(completionMask_10_reset),
    .io_in(completionMask_10_io_in),
    .io_out(completionMask_10_io_out),
    .io_enable(completionMask_10_io_enable)
  );
  FF_9 completionMask_11 (
    .clock(completionMask_11_clock),
    .reset(completionMask_11_reset),
    .io_in(completionMask_11_io_in),
    .io_out(completionMask_11_io_out),
    .io_enable(completionMask_11_io_enable)
  );
  FF_9 completionMask_12 (
    .clock(completionMask_12_clock),
    .reset(completionMask_12_reset),
    .io_in(completionMask_12_io_in),
    .io_out(completionMask_12_io_out),
    .io_enable(completionMask_12_io_enable)
  );
  FF_9 completionMask_13 (
    .clock(completionMask_13_clock),
    .reset(completionMask_13_reset),
    .io_in(completionMask_13_io_in),
    .io_out(completionMask_13_io_out),
    .io_enable(completionMask_13_io_enable)
  );
  FF_9 completionMask_14 (
    .clock(completionMask_14_clock),
    .reset(completionMask_14_reset),
    .io_in(completionMask_14_io_in),
    .io_out(completionMask_14_io_out),
    .io_enable(completionMask_14_io_enable)
  );
  FF_9 completionMask_15 (
    .clock(completionMask_15_clock),
    .reset(completionMask_15_reset),
    .io_in(completionMask_15_io_in),
    .io_out(completionMask_15_io_out),
    .io_enable(completionMask_15_io_enable)
  );
  SRFF_sp wasSparseWren (
    .clock(wasSparseWren_clock),
    .reset(wasSparseWren_reset),
    .io_input_set(wasSparseWren_io_input_set),
    .io_input_reset(wasSparseWren_io_input_reset),
    .io_input_asyn_reset(wasSparseWren_io_input_asyn_reset),
    .io_output_data(wasSparseWren_io_output_data)
  );
  WidthConverterFIFO rdataFifos_0 (
    .clock(rdataFifos_0_clock),
    .reset(rdataFifos_0_reset),
    .io_enqVld(rdataFifos_0_io_enqVld),
    .io_full(rdataFifos_0_io_full),
    .io_empty(rdataFifos_0_io_empty),
    .io_almostFull(rdataFifos_0_io_almostFull)
  );
  FIFOCounter wrespFifos_0 (
    .clock(wrespFifos_0_clock),
    .reset(wrespFifos_0_reset),
    .io_enqVld(wrespFifos_0_io_enqVld),
    .io_full(wrespFifos_0_io_full),
    .io_almostFull(wrespFifos_0_io_almostFull)
  );
  MuxNType_17 MuxNType_1 (
    .io_ins_0(MuxNType_1_io_ins_0),
    .io_out(MuxNType_1_io_out)
  );
  MuxNType_17 MuxNType_2 (
    .io_ins_0(MuxNType_2_io_ins_0),
    .io_out(MuxNType_2_io_out)
  );
  Counter_19 Counter (
    .clock(Counter_clock),
    .reset(Counter_reset),
    .io_max(Counter_io_max),
    .io_out(Counter_io_out),
    .io_enable(Counter_io_enable),
    .io_saturate(Counter_io_saturate),
    .io_done(Counter_io_done)
  );
  Counter_12 Counter_1 (
    .clock(Counter_1_clock),
    .reset(Counter_1_reset),
    .io_max(Counter_1_io_max),
    .io_out(Counter_1_io_out),
    .io_enable(Counter_1_io_enable),
    .io_done(Counter_1_io_done)
  );
  FF_42 FF (
    .clock(FF_clock),
    .reset(FF_reset),
    .io_in(FF_io_in),
    .io_init(FF_io_init),
    .io_out(FF_io_out),
    .io_enable(FF_io_enable)
  );
  FF_42 FF_1 (
    .clock(FF_1_clock),
    .reset(FF_1_reset),
    .io_in(FF_1_io_in),
    .io_init(FF_1_io_init),
    .io_out(FF_1_io_out),
    .io_enable(FF_1_io_enable)
  );
  FF_42 FF_2 (
    .clock(FF_2_clock),
    .reset(FF_2_reset),
    .io_in(FF_2_io_in),
    .io_init(FF_2_io_init),
    .io_out(FF_2_io_out),
    .io_enable(FF_2_io_enable)
  );
  FF_42 FF_3 (
    .clock(FF_3_clock),
    .reset(FF_3_reset),
    .io_in(FF_3_io_in),
    .io_init(FF_3_io_init),
    .io_out(FF_3_io_out),
    .io_enable(FF_3_io_enable)
  );
  FF_42 FF_4 (
    .clock(FF_4_clock),
    .reset(FF_4_reset),
    .io_in(FF_4_io_in),
    .io_init(FF_4_io_init),
    .io_out(FF_4_io_out),
    .io_enable(FF_4_io_enable)
  );
  FF_42 FF_5 (
    .clock(FF_5_clock),
    .reset(FF_5_reset),
    .io_in(FF_5_io_in),
    .io_init(FF_5_io_init),
    .io_out(FF_5_io_out),
    .io_enable(FF_5_io_enable)
  );
  FF_42 FF_6 (
    .clock(FF_6_clock),
    .reset(FF_6_reset),
    .io_in(FF_6_io_in),
    .io_init(FF_6_io_init),
    .io_out(FF_6_io_out),
    .io_enable(FF_6_io_enable)
  );
  FF_42 FF_7 (
    .clock(FF_7_clock),
    .reset(FF_7_reset),
    .io_in(FF_7_io_in),
    .io_init(FF_7_io_init),
    .io_out(FF_7_io_out),
    .io_enable(FF_7_io_enable)
  );
  FF_42 FF_8 (
    .clock(FF_8_clock),
    .reset(FF_8_reset),
    .io_in(FF_8_io_in),
    .io_init(FF_8_io_init),
    .io_out(FF_8_io_out),
    .io_enable(FF_8_io_enable)
  );
  FF_42 FF_9 (
    .clock(FF_9_clock),
    .reset(FF_9_reset),
    .io_in(FF_9_io_in),
    .io_init(FF_9_io_init),
    .io_out(FF_9_io_out),
    .io_enable(FF_9_io_enable)
  );
  FF_42 FF_10 (
    .clock(FF_10_clock),
    .reset(FF_10_reset),
    .io_in(FF_10_io_in),
    .io_init(FF_10_io_init),
    .io_out(FF_10_io_out),
    .io_enable(FF_10_io_enable)
  );
  FF_42 FF_11 (
    .clock(FF_11_clock),
    .reset(FF_11_reset),
    .io_in(FF_11_io_in),
    .io_init(FF_11_io_init),
    .io_out(FF_11_io_out),
    .io_enable(FF_11_io_enable)
  );
  FF_42 FF_12 (
    .clock(FF_12_clock),
    .reset(FF_12_reset),
    .io_in(FF_12_io_in),
    .io_init(FF_12_io_init),
    .io_out(FF_12_io_out),
    .io_enable(FF_12_io_enable)
  );
  FF_42 FF_13 (
    .clock(FF_13_clock),
    .reset(FF_13_reset),
    .io_in(FF_13_io_in),
    .io_init(FF_13_io_init),
    .io_out(FF_13_io_out),
    .io_enable(FF_13_io_enable)
  );
  FF_42 FF_14 (
    .clock(FF_14_clock),
    .reset(FF_14_reset),
    .io_in(FF_14_io_in),
    .io_init(FF_14_io_init),
    .io_out(FF_14_io_out),
    .io_enable(FF_14_io_enable)
  );
  FF_42 FF_15 (
    .clock(FF_15_clock),
    .reset(FF_15_reset),
    .io_in(FF_15_io_in),
    .io_init(FF_15_io_init),
    .io_out(FF_15_io_out),
    .io_enable(FF_15_io_enable)
  );
  FF_42 FF_16 (
    .clock(FF_16_clock),
    .reset(FF_16_reset),
    .io_in(FF_16_io_in),
    .io_init(FF_16_io_init),
    .io_out(FF_16_io_out),
    .io_enable(FF_16_io_enable)
  );
  FF_42 FF_17 (
    .clock(FF_17_clock),
    .reset(FF_17_reset),
    .io_in(FF_17_io_in),
    .io_init(FF_17_io_init),
    .io_out(FF_17_io_out),
    .io_enable(FF_17_io_enable)
  );
  FF_42 FF_18 (
    .clock(FF_18_clock),
    .reset(FF_18_reset),
    .io_in(FF_18_io_in),
    .io_init(FF_18_io_init),
    .io_out(FF_18_io_out),
    .io_enable(FF_18_io_enable)
  );
  FF_42 FF_19 (
    .clock(FF_19_clock),
    .reset(FF_19_reset),
    .io_in(FF_19_io_in),
    .io_init(FF_19_io_init),
    .io_out(FF_19_io_out),
    .io_enable(FF_19_io_enable)
  );
  FF_42 FF_20 (
    .clock(FF_20_clock),
    .reset(FF_20_reset),
    .io_in(FF_20_io_in),
    .io_init(FF_20_io_init),
    .io_out(FF_20_io_out),
    .io_enable(FF_20_io_enable)
  );
  FF_42 FF_21 (
    .clock(FF_21_clock),
    .reset(FF_21_reset),
    .io_in(FF_21_io_in),
    .io_init(FF_21_io_init),
    .io_out(FF_21_io_out),
    .io_enable(FF_21_io_enable)
  );
  FF_42 FF_22 (
    .clock(FF_22_clock),
    .reset(FF_22_reset),
    .io_in(FF_22_io_in),
    .io_init(FF_22_io_init),
    .io_out(FF_22_io_out),
    .io_enable(FF_22_io_enable)
  );
  FF_42 FF_23 (
    .clock(FF_23_clock),
    .reset(FF_23_reset),
    .io_in(FF_23_io_in),
    .io_init(FF_23_io_init),
    .io_out(FF_23_io_out),
    .io_enable(FF_23_io_enable)
  );
  FF_42 FF_24 (
    .clock(FF_24_clock),
    .reset(FF_24_reset),
    .io_in(FF_24_io_in),
    .io_init(FF_24_io_init),
    .io_out(FF_24_io_out),
    .io_enable(FF_24_io_enable)
  );
  FF_42 FF_25 (
    .clock(FF_25_clock),
    .reset(FF_25_reset),
    .io_in(FF_25_io_in),
    .io_init(FF_25_io_init),
    .io_out(FF_25_io_out),
    .io_enable(FF_25_io_enable)
  );
  FF_42 FF_26 (
    .clock(FF_26_clock),
    .reset(FF_26_reset),
    .io_in(FF_26_io_in),
    .io_init(FF_26_io_init),
    .io_out(FF_26_io_out),
    .io_enable(FF_26_io_enable)
  );
  FF_42 FF_27 (
    .clock(FF_27_clock),
    .reset(FF_27_reset),
    .io_in(FF_27_io_in),
    .io_init(FF_27_io_init),
    .io_out(FF_27_io_out),
    .io_enable(FF_27_io_enable)
  );
  FF_42 FF_28 (
    .clock(FF_28_clock),
    .reset(FF_28_reset),
    .io_in(FF_28_io_in),
    .io_init(FF_28_io_init),
    .io_out(FF_28_io_out),
    .io_enable(FF_28_io_enable)
  );
  FF_42 FF_29 (
    .clock(FF_29_clock),
    .reset(FF_29_reset),
    .io_in(FF_29_io_in),
    .io_init(FF_29_io_init),
    .io_out(FF_29_io_out),
    .io_enable(FF_29_io_enable)
  );
  FF_42 FF_30 (
    .clock(FF_30_clock),
    .reset(FF_30_reset),
    .io_in(FF_30_io_in),
    .io_init(FF_30_io_init),
    .io_out(FF_30_io_out),
    .io_enable(FF_30_io_enable)
  );
  FF_42 FF_31 (
    .clock(FF_31_clock),
    .reset(FF_31_reset),
    .io_in(FF_31_io_in),
    .io_init(FF_31_io_init),
    .io_out(FF_31_io_out),
    .io_enable(FF_31_io_enable)
  );
  Counter_12 Counter_2 (
    .clock(Counter_2_clock),
    .reset(Counter_2_reset),
    .io_max(Counter_2_io_max),
    .io_out(Counter_2_io_out),
    .io_enable(Counter_2_io_enable),
    .io_done(Counter_2_io_done)
  );
  Counter_12 Counter_3 (
    .clock(Counter_3_clock),
    .reset(Counter_3_reset),
    .io_max(Counter_3_io_max),
    .io_out(Counter_3_io_out),
    .io_enable(Counter_3_io_enable),
    .io_done(Counter_3_io_done)
  );
  Counter_12 Counter_4 (
    .clock(Counter_4_clock),
    .reset(Counter_4_reset),
    .io_max(Counter_4_io_max),
    .io_out(Counter_4_io_out),
    .io_enable(Counter_4_io_enable),
    .io_done(Counter_4_io_done)
  );
  Counter_12 Counter_5 (
    .clock(Counter_5_clock),
    .reset(Counter_5_reset),
    .io_max(Counter_5_io_max),
    .io_out(Counter_5_io_out),
    .io_enable(Counter_5_io_enable),
    .io_done(Counter_5_io_done)
  );
  Counter_12 Counter_6 (
    .clock(Counter_6_clock),
    .reset(Counter_6_reset),
    .io_max(Counter_6_io_max),
    .io_out(Counter_6_io_out),
    .io_enable(Counter_6_io_enable),
    .io_done(Counter_6_io_done)
  );
  Counter_12 Counter_7 (
    .clock(Counter_7_clock),
    .reset(Counter_7_reset),
    .io_max(Counter_7_io_max),
    .io_out(Counter_7_io_out),
    .io_enable(Counter_7_io_enable),
    .io_done(Counter_7_io_done)
  );
  Counter_12 Counter_8 (
    .clock(Counter_8_clock),
    .reset(Counter_8_reset),
    .io_max(Counter_8_io_max),
    .io_out(Counter_8_io_out),
    .io_enable(Counter_8_io_enable),
    .io_done(Counter_8_io_done)
  );
  Counter_12 Counter_9 (
    .clock(Counter_9_clock),
    .reset(Counter_9_reset),
    .io_max(Counter_9_io_max),
    .io_out(Counter_9_io_out),
    .io_enable(Counter_9_io_enable),
    .io_done(Counter_9_io_done)
  );
  Counter_12 Counter_10 (
    .clock(Counter_10_clock),
    .reset(Counter_10_reset),
    .io_max(Counter_10_io_max),
    .io_out(Counter_10_io_out),
    .io_enable(Counter_10_io_enable),
    .io_done(Counter_10_io_done)
  );
  Counter_12 Counter_11 (
    .clock(Counter_11_clock),
    .reset(Counter_11_reset),
    .io_max(Counter_11_io_max),
    .io_out(Counter_11_io_out),
    .io_enable(Counter_11_io_enable),
    .io_done(Counter_11_io_done)
  );
  Counter_12 Counter_12 (
    .clock(Counter_12_clock),
    .reset(Counter_12_reset),
    .io_max(Counter_12_io_max),
    .io_out(Counter_12_io_out),
    .io_enable(Counter_12_io_enable),
    .io_done(Counter_12_io_done)
  );
  Counter_12 Counter_13 (
    .clock(Counter_13_clock),
    .reset(Counter_13_reset),
    .io_max(Counter_13_io_max),
    .io_out(Counter_13_io_out),
    .io_enable(Counter_13_io_enable),
    .io_done(Counter_13_io_done)
  );
  FF_1160 FF_32 (
    .clock(FF_32_clock),
    .reset(FF_32_reset),
    .io_in(FF_32_io_in),
    .io_init(FF_32_io_init),
    .io_out(FF_32_io_out),
    .io_enable(FF_32_io_enable)
  );
  FF_1160 FF_33 (
    .clock(FF_33_clock),
    .reset(FF_33_reset),
    .io_in(FF_33_io_in),
    .io_init(FF_33_io_init),
    .io_out(FF_33_io_out),
    .io_enable(FF_33_io_enable)
  );
  Counter_12 Counter_14 (
    .clock(Counter_14_clock),
    .reset(Counter_14_reset),
    .io_max(Counter_14_io_max),
    .io_out(Counter_14_io_out),
    .io_enable(Counter_14_io_enable),
    .io_done(Counter_14_io_done)
  );
  Counter_12 Counter_15 (
    .clock(Counter_15_clock),
    .reset(Counter_15_reset),
    .io_max(Counter_15_io_max),
    .io_out(Counter_15_io_out),
    .io_enable(Counter_15_io_enable),
    .io_done(Counter_15_io_done)
  );
  Counter_12 Counter_16 (
    .clock(Counter_16_clock),
    .reset(Counter_16_reset),
    .io_max(Counter_16_io_max),
    .io_out(Counter_16_io_out),
    .io_enable(Counter_16_io_enable),
    .io_done(Counter_16_io_done)
  );
  Counter_12 Counter_17 (
    .clock(Counter_17_clock),
    .reset(Counter_17_reset),
    .io_max(Counter_17_io_max),
    .io_out(Counter_17_io_out),
    .io_enable(Counter_17_io_enable),
    .io_done(Counter_17_io_done)
  );
  Counter_12 Counter_18 (
    .clock(Counter_18_clock),
    .reset(Counter_18_reset),
    .io_max(Counter_18_io_max),
    .io_out(Counter_18_io_out),
    .io_enable(Counter_18_io_enable),
    .io_done(Counter_18_io_done)
  );
  Counter_12 Counter_19 (
    .clock(Counter_19_clock),
    .reset(Counter_19_reset),
    .io_max(Counter_19_io_max),
    .io_out(Counter_19_io_out),
    .io_enable(Counter_19_io_enable),
    .io_done(Counter_19_io_done)
  );
  Counter_12 Counter_20 (
    .clock(Counter_20_clock),
    .reset(Counter_20_reset),
    .io_max(Counter_20_io_max),
    .io_out(Counter_20_io_out),
    .io_enable(Counter_20_io_enable),
    .io_done(Counter_20_io_done)
  );
  Counter_12 Counter_21 (
    .clock(Counter_21_clock),
    .reset(Counter_21_reset),
    .io_max(Counter_21_io_max),
    .io_out(Counter_21_io_out),
    .io_enable(Counter_21_io_enable),
    .io_done(Counter_21_io_done)
  );
  Counter_12 Counter_22 (
    .clock(Counter_22_clock),
    .reset(Counter_22_reset),
    .io_max(Counter_22_io_max),
    .io_out(Counter_22_io_out),
    .io_enable(Counter_22_io_enable),
    .io_done(Counter_22_io_done)
  );
  Counter_12 Counter_23 (
    .clock(Counter_23_clock),
    .reset(Counter_23_reset),
    .io_max(Counter_23_io_max),
    .io_out(Counter_23_io_out),
    .io_enable(Counter_23_io_enable),
    .io_done(Counter_23_io_done)
  );
  Counter_12 Counter_24 (
    .clock(Counter_24_clock),
    .reset(Counter_24_reset),
    .io_max(Counter_24_io_max),
    .io_out(Counter_24_io_out),
    .io_enable(Counter_24_io_enable),
    .io_done(Counter_24_io_done)
  );
  Counter_12 Counter_25 (
    .clock(Counter_25_clock),
    .reset(Counter_25_reset),
    .io_max(Counter_25_io_max),
    .io_out(Counter_25_io_out),
    .io_enable(Counter_25_io_enable),
    .io_done(Counter_25_io_done)
  );
  Counter_12 Counter_26 (
    .clock(Counter_26_clock),
    .reset(Counter_26_reset),
    .io_max(Counter_26_io_max),
    .io_out(Counter_26_io_out),
    .io_enable(Counter_26_io_enable),
    .io_done(Counter_26_io_done)
  );
  assign _T_485 = commandFifo_io_deq_0[81:18];
  assign _T_486 = commandFifo_io_deq_0[17];
  assign _T_487 = commandFifo_io_deq_0[16];
  assign _T_488 = commandFifo_io_deq_0[15:0];
  assign _T_495 = ~ commandFifo_io_empty;
  assign isSparse = headCommand_isSparse & _T_495;
  assign _T_497 = headCommand_size[15:6];
  assign _T_498 = headCommand_size[5:0];
  assign _T_500 = _T_498 != 6'h0;
  assign _GEN_0 = {{9'd0}, _T_500};
  assign _T_501 = _T_497 + _GEN_0;
  assign sizeInBursts = _T_501[9:0];
  assign _T_506 = wrPhase_io_output_data | headCommand_isWr;
  assign writeCmd = _T_495 & _T_506;
  assign _T_507 = ~ wdataFifo_io_empty;
  assign wdataValid = writeCmd & _T_507;
  assign _T_509 = commandFifo_io_tag - 1'h1;
  assign _T_510 = $unsigned(_T_509);
  assign _T_511 = _T_510[0:0];
  assign _T_513 = commandFifo_io_tag >= 1'h1;
  assign _T_515 = isSparse & headCommand_isWr;
  assign _T_517 = _T_515 & _T_495;
  assign _T_525 = writeCmd ? sizeInBursts : 10'h1;
  assign _T_536 = burstVld & headCommand_isWr;
  assign _T_537 = burstCounter_io_done | _T_536;
  assign _T_540 = burstCounter_io_done ? 1'h0 : dramReadySeen;
  assign _T_544 = io_enable & _T_495;
  assign _T_545 = ~ dramReadySeen;
  assign _T_546 = wdataValid & _T_545;
  assign _T_548 = writeCmd ? _T_546 : 1'h1;
  assign _T_549 = _T_544 & _T_548;
  assign elementID = burstTagCounter_io_out[3:0];
  assign _T_567 = ~ _T_515;
  assign _T_580 = burstCounter_io_done;
  assign validMask_0 = ccache_io_rmetaData_0[4];
  assign validMask_1 = ccache_io_rmetaData_1[4];
  assign validMask_2 = ccache_io_rmetaData_2[4];
  assign validMask_3 = ccache_io_rmetaData_3[4];
  assign validMask_4 = ccache_io_rmetaData_4[4];
  assign validMask_5 = ccache_io_rmetaData_5[4];
  assign validMask_6 = ccache_io_rmetaData_6[4];
  assign validMask_7 = ccache_io_rmetaData_7[4];
  assign validMask_8 = ccache_io_rmetaData_8[4];
  assign validMask_9 = ccache_io_rmetaData_9[4];
  assign validMask_10 = ccache_io_rmetaData_10[4];
  assign validMask_11 = ccache_io_rmetaData_11[4];
  assign validMask_12 = ccache_io_rmetaData_12[4];
  assign validMask_13 = ccache_io_rmetaData_13[4];
  assign validMask_14 = ccache_io_rmetaData_14[4];
  assign validMask_15 = ccache_io_rmetaData_15[4];
  assign _T_845 = sizeInBursts - 10'h1;
  assign _T_846 = $unsigned(_T_845);
  assign _T_847 = _T_846[9:0];
  assign _GEN_1 = {{22'd0}, _T_847};
  assign _T_848 = burstCounter_io_out == _GEN_1;
  assign wlast = wdataValid & _T_848;
  assign _T_849 = ~ sparseWriteEnable;
  assign _T_852 = _T_495 & headCommand_isWr;
  assign _T_853 = wlast | wasSparseWren_io_output_data;
  assign _T_869 = rdataFifos_0_io_full | rdataFifos_0_io_almostFull;
  assign _T_870 = ~ _T_869;
  assign _T_890 = wrespFifos_0_io_full | wrespFifos_0_io_almostFull;
  assign _T_891 = ~ _T_890;
  assign _T_1241 = ~ io_dram_rresp_ready;
  assign _T_1249 = io_enable & io_dram_rresp_ready;
  assign _T_1257 = io_enable & _T_1241;
  assign io_debugSignals_0 = Counter_io_out[31:0];
  assign io_debugSignals_1 = FF_io_out;
  assign io_debugSignals_2 = FF_1_io_out;
  assign io_debugSignals_3 = FF_2_io_out;
  assign io_debugSignals_4 = FF_3_io_out;
  assign io_debugSignals_5 = FF_4_io_out;
  assign io_debugSignals_6 = FF_5_io_out;
  assign io_debugSignals_7 = FF_6_io_out;
  assign io_debugSignals_8 = FF_7_io_out;
  assign io_debugSignals_9 = FF_8_io_out;
  assign io_debugSignals_10 = FF_9_io_out;
  assign io_debugSignals_11 = FF_10_io_out;
  assign io_debugSignals_12 = FF_11_io_out;
  assign io_debugSignals_13 = FF_12_io_out;
  assign io_debugSignals_14 = FF_13_io_out;
  assign io_debugSignals_15 = FF_14_io_out;
  assign io_debugSignals_16 = FF_15_io_out;
  assign io_debugSignals_17 = FF_16_io_out;
  assign io_debugSignals_18 = FF_17_io_out;
  assign io_debugSignals_19 = FF_18_io_out;
  assign io_debugSignals_20 = FF_19_io_out;
  assign io_debugSignals_21 = FF_20_io_out;
  assign io_debugSignals_22 = FF_21_io_out;
  assign io_debugSignals_23 = FF_22_io_out;
  assign io_debugSignals_24 = FF_23_io_out;
  assign io_debugSignals_25 = FF_24_io_out;
  assign io_debugSignals_26 = FF_25_io_out;
  assign io_debugSignals_27 = FF_26_io_out;
  assign io_debugSignals_28 = FF_27_io_out;
  assign io_debugSignals_29 = FF_28_io_out;
  assign io_debugSignals_30 = FF_29_io_out;
  assign io_debugSignals_31 = FF_30_io_out;
  assign io_debugSignals_32 = FF_31_io_out;
  assign io_debugSignals_33 = Counter_4_io_out;
  assign io_debugSignals_34 = Counter_5_io_out;
  assign io_debugSignals_35 = Counter_6_io_out;
  assign io_debugSignals_36 = Counter_7_io_out;
  assign io_debugSignals_37 = Counter_8_io_out;
  assign io_debugSignals_38 = Counter_9_io_out;
  assign io_debugSignals_39 = Counter_10_io_out;
  assign io_debugSignals_40 = Counter_11_io_out;
  assign io_debugSignals_41 = Counter_12_io_out;
  assign io_debugSignals_42 = Counter_13_io_out;
  assign io_debugSignals_43 = FF_33_io_out[31:0];
  assign io_debugSignals_44 = FF_32_io_out[31:0];
  assign io_debugSignals_45 = Counter_14_io_out;
  assign io_debugSignals_46 = Counter_15_io_out;
  assign io_debugSignals_47 = Counter_16_io_out;
  assign io_debugSignals_48 = Counter_17_io_out;
  assign io_debugSignals_49 = Counter_18_io_out;
  assign io_debugSignals_50 = Counter_19_io_out;
  assign io_debugSignals_51 = Counter_20_io_out;
  assign io_debugSignals_52 = Counter_21_io_out;
  assign io_debugSignals_53 = Counter_22_io_out;
  assign io_debugSignals_54 = Counter_23_io_out;
  assign io_debugSignals_55 = Counter_24_io_out;
  assign io_debugSignals_56 = Counter_25_io_out;
  assign io_debugSignals_57 = Counter_26_io_out;
  assign io_debugSignals_58 = Counter_2_io_out;
  assign io_dram_rresp_ready = MuxNType_1_io_out;
  assign commandFifo_io_deqVld = _T_580;
  assign commandFifo_clock = clock;
  assign commandFifo_reset = reset;
  assign headCommand_addr = _T_484_addr;
  assign headCommand_isWr = _T_484_isWr;
  assign headCommand_isSparse = _T_484_isSparse;
  assign headCommand_size = _T_484_size;
  assign _T_484_addr = _T_485;
  assign _T_484_isWr = _T_486;
  assign _T_484_isSparse = _T_487;
  assign _T_484_size = _T_488;
  assign wdataFifo_io_forceTag_valid = _T_513;
  assign wdataFifo_io_forceTag_bits = _T_511;
  assign wdataFifo_clock = clock;
  assign wdataFifo_reset = reset;
  assign wrPhase_io_input_set = _T_852;
  assign wrPhase_io_input_reset = _T_856;
  assign wrPhase_io_input_asyn_reset = 1'h0;
  assign wrPhase_clock = clock;
  assign wrPhase_reset = reset;
  assign burstVld = _T_549;
  assign sparseWriteEnable = _T_517;
  assign issuedFF_io_in = 1'h0;
  assign issuedFF_io_enable = 1'h1;
  assign issuedFF_clock = clock;
  assign issuedFF_reset = reset;
  assign burstCounter_io_max = {{22'd0}, _T_525};
  assign burstCounter_io_enable = 1'h0;
  assign burstCounter_clock = clock;
  assign burstCounter_reset = reset;
  assign dramReadySeen = dramReadyFF_io_out;
  assign dramReadyFF_io_in = _T_540;
  assign dramReadyFF_io_enable = _T_537;
  assign dramReadyFF_clock = clock;
  assign dramReadyFF_reset = reset;
  assign burstTagCounter_clock = clock;
  assign burstTagCounter_reset = reset;
  assign wdataSelectCounter_io_reset = _T_567;
  assign wdataSelectCounter_clock = clock;
  assign wdataSelectCounter_reset = reset;
  assign ccache_io_waddr = headCommand_addr[31:0];
  assign ccache_io_position = elementID;
  assign ccache_clock = clock;
  assign ccache_reset = reset;
  assign sgValidDepulser_io_in = 1'h0;
  assign sgValidDepulser_io_rst = 1'h0;
  assign sgValidDepulser_clock = clock;
  assign sgValidDepulser_reset = reset;
  assign gatherBuffer_0_io_in = 32'h0;
  assign gatherBuffer_0_io_init = 32'h0;
  assign gatherBuffer_0_io_enable = 1'h0;
  assign gatherBuffer_0_clock = clock;
  assign gatherBuffer_0_reset = reset;
  assign gatherBuffer_1_io_in = 32'h0;
  assign gatherBuffer_1_io_init = 32'h0;
  assign gatherBuffer_1_io_enable = 1'h0;
  assign gatherBuffer_1_clock = clock;
  assign gatherBuffer_1_reset = reset;
  assign gatherBuffer_2_io_in = 32'h0;
  assign gatherBuffer_2_io_init = 32'h0;
  assign gatherBuffer_2_io_enable = 1'h0;
  assign gatherBuffer_2_clock = clock;
  assign gatherBuffer_2_reset = reset;
  assign gatherBuffer_3_io_in = 32'h0;
  assign gatherBuffer_3_io_init = 32'h0;
  assign gatherBuffer_3_io_enable = 1'h0;
  assign gatherBuffer_3_clock = clock;
  assign gatherBuffer_3_reset = reset;
  assign gatherBuffer_4_io_in = 32'h0;
  assign gatherBuffer_4_io_init = 32'h0;
  assign gatherBuffer_4_io_enable = 1'h0;
  assign gatherBuffer_4_clock = clock;
  assign gatherBuffer_4_reset = reset;
  assign gatherBuffer_5_io_in = 32'h0;
  assign gatherBuffer_5_io_init = 32'h0;
  assign gatherBuffer_5_io_enable = 1'h0;
  assign gatherBuffer_5_clock = clock;
  assign gatherBuffer_5_reset = reset;
  assign gatherBuffer_6_io_in = 32'h0;
  assign gatherBuffer_6_io_init = 32'h0;
  assign gatherBuffer_6_io_enable = 1'h0;
  assign gatherBuffer_6_clock = clock;
  assign gatherBuffer_6_reset = reset;
  assign gatherBuffer_7_io_in = 32'h0;
  assign gatherBuffer_7_io_init = 32'h0;
  assign gatherBuffer_7_io_enable = 1'h0;
  assign gatherBuffer_7_clock = clock;
  assign gatherBuffer_7_reset = reset;
  assign gatherBuffer_8_io_in = 32'h0;
  assign gatherBuffer_8_io_init = 32'h0;
  assign gatherBuffer_8_io_enable = 1'h0;
  assign gatherBuffer_8_clock = clock;
  assign gatherBuffer_8_reset = reset;
  assign gatherBuffer_9_io_in = 32'h0;
  assign gatherBuffer_9_io_init = 32'h0;
  assign gatherBuffer_9_io_enable = 1'h0;
  assign gatherBuffer_9_clock = clock;
  assign gatherBuffer_9_reset = reset;
  assign gatherBuffer_10_io_in = 32'h0;
  assign gatherBuffer_10_io_init = 32'h0;
  assign gatherBuffer_10_io_enable = 1'h0;
  assign gatherBuffer_10_clock = clock;
  assign gatherBuffer_10_reset = reset;
  assign gatherBuffer_11_io_in = 32'h0;
  assign gatherBuffer_11_io_init = 32'h0;
  assign gatherBuffer_11_io_enable = 1'h0;
  assign gatherBuffer_11_clock = clock;
  assign gatherBuffer_11_reset = reset;
  assign gatherBuffer_12_io_in = 32'h0;
  assign gatherBuffer_12_io_init = 32'h0;
  assign gatherBuffer_12_io_enable = 1'h0;
  assign gatherBuffer_12_clock = clock;
  assign gatherBuffer_12_reset = reset;
  assign gatherBuffer_13_io_in = 32'h0;
  assign gatherBuffer_13_io_init = 32'h0;
  assign gatherBuffer_13_io_enable = 1'h0;
  assign gatherBuffer_13_clock = clock;
  assign gatherBuffer_13_reset = reset;
  assign gatherBuffer_14_io_in = 32'h0;
  assign gatherBuffer_14_io_init = 32'h0;
  assign gatherBuffer_14_io_enable = 1'h0;
  assign gatherBuffer_14_clock = clock;
  assign gatherBuffer_14_reset = reset;
  assign gatherBuffer_15_io_in = 32'h0;
  assign gatherBuffer_15_io_init = 32'h0;
  assign gatherBuffer_15_io_enable = 1'h0;
  assign gatherBuffer_15_clock = clock;
  assign gatherBuffer_15_reset = reset;
  assign completionMask_0_io_in = validMask_0;
  assign completionMask_0_io_enable = 1'h0;
  assign completionMask_0_clock = clock;
  assign completionMask_0_reset = reset;
  assign completionMask_1_io_in = validMask_1;
  assign completionMask_1_io_enable = 1'h0;
  assign completionMask_1_clock = clock;
  assign completionMask_1_reset = reset;
  assign completionMask_2_io_in = validMask_2;
  assign completionMask_2_io_enable = 1'h0;
  assign completionMask_2_clock = clock;
  assign completionMask_2_reset = reset;
  assign completionMask_3_io_in = validMask_3;
  assign completionMask_3_io_enable = 1'h0;
  assign completionMask_3_clock = clock;
  assign completionMask_3_reset = reset;
  assign completionMask_4_io_in = validMask_4;
  assign completionMask_4_io_enable = 1'h0;
  assign completionMask_4_clock = clock;
  assign completionMask_4_reset = reset;
  assign completionMask_5_io_in = validMask_5;
  assign completionMask_5_io_enable = 1'h0;
  assign completionMask_5_clock = clock;
  assign completionMask_5_reset = reset;
  assign completionMask_6_io_in = validMask_6;
  assign completionMask_6_io_enable = 1'h0;
  assign completionMask_6_clock = clock;
  assign completionMask_6_reset = reset;
  assign completionMask_7_io_in = validMask_7;
  assign completionMask_7_io_enable = 1'h0;
  assign completionMask_7_clock = clock;
  assign completionMask_7_reset = reset;
  assign completionMask_8_io_in = validMask_8;
  assign completionMask_8_io_enable = 1'h0;
  assign completionMask_8_clock = clock;
  assign completionMask_8_reset = reset;
  assign completionMask_9_io_in = validMask_9;
  assign completionMask_9_io_enable = 1'h0;
  assign completionMask_9_clock = clock;
  assign completionMask_9_reset = reset;
  assign completionMask_10_io_in = validMask_10;
  assign completionMask_10_io_enable = 1'h0;
  assign completionMask_10_clock = clock;
  assign completionMask_10_reset = reset;
  assign completionMask_11_io_in = validMask_11;
  assign completionMask_11_io_enable = 1'h0;
  assign completionMask_11_clock = clock;
  assign completionMask_11_reset = reset;
  assign completionMask_12_io_in = validMask_12;
  assign completionMask_12_io_enable = 1'h0;
  assign completionMask_12_clock = clock;
  assign completionMask_12_reset = reset;
  assign completionMask_13_io_in = validMask_13;
  assign completionMask_13_io_enable = 1'h0;
  assign completionMask_13_clock = clock;
  assign completionMask_13_reset = reset;
  assign completionMask_14_io_in = validMask_14;
  assign completionMask_14_io_enable = 1'h0;
  assign completionMask_14_clock = clock;
  assign completionMask_14_reset = reset;
  assign completionMask_15_io_in = validMask_15;
  assign completionMask_15_io_enable = 1'h0;
  assign completionMask_15_clock = clock;
  assign completionMask_15_reset = reset;
  assign wasSparseWren_io_input_set = sparseWriteEnable;
  assign wasSparseWren_io_input_reset = _T_849;
  assign wasSparseWren_io_input_asyn_reset = 1'h0;
  assign wasSparseWren_clock = clock;
  assign wasSparseWren_reset = reset;
  assign rdataFifos_0_io_enqVld = 1'h0;
  assign rdataFifos_0_clock = clock;
  assign rdataFifos_0_reset = reset;
  assign wrespFifos_0_io_enqVld = 1'h0;
  assign wrespFifos_0_clock = clock;
  assign wrespFifos_0_reset = reset;
  assign MuxNType_1_io_ins_0 = _T_886_0;
  assign _T_886_0 = _T_870;
  assign MuxNType_2_io_ins_0 = _T_894_0;
  assign _T_894_0 = _T_891;
  assign Counter_io_max = 40'hffffffffff;
  assign Counter_io_enable = io_enable;
  assign Counter_io_saturate = 1'h0;
  assign Counter_clock = clock;
  assign Counter_reset = reset;
  assign Counter_1_io_max = 32'hffffffff;
  assign Counter_1_io_enable = 1'h0;
  assign Counter_1_clock = clock;
  assign Counter_1_reset = reset;
  assign FF_io_in = 32'h0;
  assign FF_io_init = 32'h175bf;
  assign FF_io_enable = 1'h0;
  assign FF_clock = clock;
  assign FF_reset = reset;
  assign FF_1_io_in = 32'h0;
  assign FF_1_io_init = 32'h2eb7e;
  assign FF_1_io_enable = 1'h0;
  assign FF_1_clock = clock;
  assign FF_1_reset = reset;
  assign FF_2_io_in = 32'h0;
  assign FF_2_io_init = 32'h2eb7f;
  assign FF_2_io_enable = 1'h0;
  assign FF_2_clock = clock;
  assign FF_2_reset = reset;
  assign FF_3_io_in = 32'h0;
  assign FF_3_io_init = 32'h5d6fc;
  assign FF_3_io_enable = 1'h0;
  assign FF_3_clock = clock;
  assign FF_3_reset = reset;
  assign FF_4_io_in = 32'h0;
  assign FF_4_io_init = 32'h5d6fd;
  assign FF_4_io_enable = 1'h0;
  assign FF_4_clock = clock;
  assign FF_4_reset = reset;
  assign FF_5_io_in = 32'h0;
  assign FF_5_io_init = 32'h5d6fe;
  assign FF_5_io_enable = 1'h0;
  assign FF_5_clock = clock;
  assign FF_5_reset = reset;
  assign FF_6_io_in = 32'h0;
  assign FF_6_io_init = 32'h5d6ff;
  assign FF_6_io_enable = 1'h0;
  assign FF_6_clock = clock;
  assign FF_6_reset = reset;
  assign FF_7_io_in = 32'h0;
  assign FF_7_io_init = 32'hbadf8;
  assign FF_7_io_enable = 1'h0;
  assign FF_7_clock = clock;
  assign FF_7_reset = reset;
  assign FF_8_io_in = 32'h0;
  assign FF_8_io_init = 32'hbadf9;
  assign FF_8_io_enable = 1'h0;
  assign FF_8_clock = clock;
  assign FF_8_reset = reset;
  assign FF_9_io_in = 32'h0;
  assign FF_9_io_init = 32'hbadfa;
  assign FF_9_io_enable = 1'h0;
  assign FF_9_clock = clock;
  assign FF_9_reset = reset;
  assign FF_10_io_in = 32'h0;
  assign FF_10_io_init = 32'hbadfb;
  assign FF_10_io_enable = 1'h0;
  assign FF_10_clock = clock;
  assign FF_10_reset = reset;
  assign FF_11_io_in = 32'h0;
  assign FF_11_io_init = 32'hbadfc;
  assign FF_11_io_enable = 1'h0;
  assign FF_11_clock = clock;
  assign FF_11_reset = reset;
  assign FF_12_io_in = 32'h0;
  assign FF_12_io_init = 32'hbadfd;
  assign FF_12_io_enable = 1'h0;
  assign FF_12_clock = clock;
  assign FF_12_reset = reset;
  assign FF_13_io_in = 32'h0;
  assign FF_13_io_init = 32'hbadfe;
  assign FF_13_io_enable = 1'h0;
  assign FF_13_clock = clock;
  assign FF_13_reset = reset;
  assign FF_14_io_in = 32'h0;
  assign FF_14_io_init = 32'hbadff;
  assign FF_14_io_enable = 1'h0;
  assign FF_14_clock = clock;
  assign FF_14_reset = reset;
  assign FF_15_io_in = 32'h0;
  assign FF_15_io_init = 32'h175bf0;
  assign FF_15_io_enable = 1'h0;
  assign FF_15_clock = clock;
  assign FF_15_reset = reset;
  assign FF_16_io_in = 32'h0;
  assign FF_16_io_init = 32'h175bf1;
  assign FF_16_io_enable = 1'h0;
  assign FF_16_clock = clock;
  assign FF_16_reset = reset;
  assign FF_17_io_in = 32'h0;
  assign FF_17_io_init = 32'h175bf2;
  assign FF_17_io_enable = 1'h0;
  assign FF_17_clock = clock;
  assign FF_17_reset = reset;
  assign FF_18_io_in = 32'h0;
  assign FF_18_io_init = 32'h175bf3;
  assign FF_18_io_enable = 1'h0;
  assign FF_18_clock = clock;
  assign FF_18_reset = reset;
  assign FF_19_io_in = 32'h0;
  assign FF_19_io_init = 32'h175bf4;
  assign FF_19_io_enable = 1'h0;
  assign FF_19_clock = clock;
  assign FF_19_reset = reset;
  assign FF_20_io_in = 32'h0;
  assign FF_20_io_init = 32'h175bf5;
  assign FF_20_io_enable = 1'h0;
  assign FF_20_clock = clock;
  assign FF_20_reset = reset;
  assign FF_21_io_in = 32'h0;
  assign FF_21_io_init = 32'h175bf6;
  assign FF_21_io_enable = 1'h0;
  assign FF_21_clock = clock;
  assign FF_21_reset = reset;
  assign FF_22_io_in = 32'h0;
  assign FF_22_io_init = 32'h175bf7;
  assign FF_22_io_enable = 1'h0;
  assign FF_22_clock = clock;
  assign FF_22_reset = reset;
  assign FF_23_io_in = 32'h0;
  assign FF_23_io_init = 32'h175bf8;
  assign FF_23_io_enable = 1'h0;
  assign FF_23_clock = clock;
  assign FF_23_reset = reset;
  assign FF_24_io_in = 32'h0;
  assign FF_24_io_init = 32'h175bf9;
  assign FF_24_io_enable = 1'h0;
  assign FF_24_clock = clock;
  assign FF_24_reset = reset;
  assign FF_25_io_in = 32'h0;
  assign FF_25_io_init = 32'h175bfa;
  assign FF_25_io_enable = 1'h0;
  assign FF_25_clock = clock;
  assign FF_25_reset = reset;
  assign FF_26_io_in = 32'h0;
  assign FF_26_io_init = 32'h175bfb;
  assign FF_26_io_enable = 1'h0;
  assign FF_26_clock = clock;
  assign FF_26_reset = reset;
  assign FF_27_io_in = 32'h0;
  assign FF_27_io_init = 32'h175bfc;
  assign FF_27_io_enable = 1'h0;
  assign FF_27_clock = clock;
  assign FF_27_reset = reset;
  assign FF_28_io_in = 32'h0;
  assign FF_28_io_init = 32'h175bfd;
  assign FF_28_io_enable = 1'h0;
  assign FF_28_clock = clock;
  assign FF_28_reset = reset;
  assign FF_29_io_in = 32'h0;
  assign FF_29_io_init = 32'h175bfe;
  assign FF_29_io_enable = 1'h0;
  assign FF_29_clock = clock;
  assign FF_29_reset = reset;
  assign FF_30_io_in = 32'h0;
  assign FF_30_io_init = 32'h175bff;
  assign FF_30_io_enable = 1'h0;
  assign FF_30_clock = clock;
  assign FF_30_reset = reset;
  assign FF_31_io_in = 32'h0;
  assign FF_31_io_init = 32'h2eb7e0;
  assign FF_31_io_enable = 1'h0;
  assign FF_31_clock = clock;
  assign FF_31_reset = reset;
  assign Counter_2_io_max = 32'hffffffff;
  assign Counter_2_io_enable = 1'h0;
  assign Counter_2_clock = clock;
  assign Counter_2_reset = reset;
  assign Counter_3_io_max = 32'hffffffff;
  assign Counter_3_io_enable = 1'h0;
  assign Counter_3_clock = clock;
  assign Counter_3_reset = reset;
  assign Counter_4_io_max = 32'hffffffff;
  assign Counter_4_io_enable = 1'h0;
  assign Counter_4_clock = clock;
  assign Counter_4_reset = reset;
  assign Counter_5_io_max = 32'hffffffff;
  assign Counter_5_io_enable = _T_544;
  assign Counter_5_clock = clock;
  assign Counter_5_reset = reset;
  assign Counter_6_io_max = 32'hffffffff;
  assign Counter_6_io_enable = 1'h0;
  assign Counter_6_clock = clock;
  assign Counter_6_reset = reset;
  assign Counter_7_io_max = 32'hffffffff;
  assign Counter_7_io_enable = 1'h0;
  assign Counter_7_clock = clock;
  assign Counter_7_reset = reset;
  assign Counter_8_io_max = 32'hffffffff;
  assign Counter_8_io_enable = 1'h0;
  assign Counter_8_clock = clock;
  assign Counter_8_reset = reset;
  assign Counter_9_io_max = 32'hffffffff;
  assign Counter_9_io_enable = 1'h0;
  assign Counter_9_clock = clock;
  assign Counter_9_reset = reset;
  assign Counter_10_io_max = 32'hffffffff;
  assign Counter_10_io_enable = 1'h0;
  assign Counter_10_clock = clock;
  assign Counter_10_reset = reset;
  assign Counter_11_io_max = 32'hffffffff;
  assign Counter_11_io_enable = 1'h0;
  assign Counter_11_clock = clock;
  assign Counter_11_reset = reset;
  assign Counter_12_io_max = 32'hffffffff;
  assign Counter_12_io_enable = 1'h0;
  assign Counter_12_clock = clock;
  assign Counter_12_reset = reset;
  assign Counter_13_io_max = 32'hffffffff;
  assign Counter_13_io_enable = 1'h0;
  assign Counter_13_clock = clock;
  assign Counter_13_reset = reset;
  assign FF_32_io_in = headCommand_addr;
  assign FF_32_io_init = 64'h2eb7e9;
  assign FF_32_io_enable = 1'h0;
  assign FF_32_clock = clock;
  assign FF_32_reset = reset;
  assign FF_33_io_in = headCommand_addr;
  assign FF_33_io_init = 64'h2eb7e9;
  assign FF_33_io_enable = 1'h1;
  assign FF_33_clock = clock;
  assign FF_33_reset = reset;
  assign Counter_14_io_max = 32'hffffffff;
  assign Counter_14_io_enable = 1'h0;
  assign Counter_14_clock = clock;
  assign Counter_14_reset = reset;
  assign Counter_15_io_max = 32'hffffffff;
  assign Counter_15_io_enable = io_enable;
  assign Counter_15_clock = clock;
  assign Counter_15_reset = reset;
  assign Counter_16_io_max = 32'hffffffff;
  assign Counter_16_io_enable = 1'h0;
  assign Counter_16_clock = clock;
  assign Counter_16_reset = reset;
  assign Counter_17_io_max = 32'hffffffff;
  assign Counter_17_io_enable = _T_1249;
  assign Counter_17_clock = clock;
  assign Counter_17_reset = reset;
  assign Counter_18_io_max = 32'hffffffff;
  assign Counter_18_io_enable = _T_1257;
  assign Counter_18_clock = clock;
  assign Counter_18_reset = reset;
  assign Counter_19_io_max = 32'hffffffff;
  assign Counter_19_io_enable = 1'h0;
  assign Counter_19_clock = clock;
  assign Counter_19_reset = reset;
  assign Counter_20_io_max = 32'hffffffff;
  assign Counter_20_io_enable = 1'h0;
  assign Counter_20_clock = clock;
  assign Counter_20_reset = reset;
  assign Counter_21_io_max = 32'hffffffff;
  assign Counter_21_io_enable = 1'h0;
  assign Counter_21_clock = clock;
  assign Counter_21_reset = reset;
  assign Counter_22_io_max = 32'hffffffff;
  assign Counter_22_io_enable = 1'h0;
  assign Counter_22_clock = clock;
  assign Counter_22_reset = reset;
  assign Counter_23_io_max = 32'hffffffff;
  assign Counter_23_io_enable = 1'h0;
  assign Counter_23_clock = clock;
  assign Counter_23_reset = reset;
  assign Counter_24_io_max = 32'hffffffff;
  assign Counter_24_io_enable = 1'h0;
  assign Counter_24_clock = clock;
  assign Counter_24_reset = reset;
  assign Counter_25_io_max = 32'hffffffff;
  assign Counter_25_io_enable = rdataFifos_0_io_enqVld;
  assign Counter_25_clock = clock;
  assign Counter_25_reset = reset;
  assign Counter_26_io_max = 32'hffffffff;
  assign Counter_26_io_enable = wrespFifos_0_io_enqVld;
  assign Counter_26_clock = clock;
  assign Counter_26_reset = reset;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  _T_856 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_856 <= 1'h0;
    end else begin
      _T_856 <= _T_853;
    end
  end
endmodule
module MuxN_6(
  input  [63:0] io_ins_0,
  input  [63:0] io_ins_1,
  input  [63:0] io_ins_2,
  input  [63:0] io_ins_3,
  input  [63:0] io_ins_4,
  input  [63:0] io_ins_5,
  input  [63:0] io_ins_6,
  input  [63:0] io_ins_7,
  input  [63:0] io_ins_8,
  input  [63:0] io_ins_9,
  input  [63:0] io_ins_10,
  input  [63:0] io_ins_11,
  input  [63:0] io_ins_12,
  input  [63:0] io_ins_13,
  input  [63:0] io_ins_14,
  input  [63:0] io_ins_15,
  input  [63:0] io_ins_16,
  input  [63:0] io_ins_17,
  input  [63:0] io_ins_18,
  input  [63:0] io_ins_19,
  input  [63:0] io_ins_20,
  input  [63:0] io_ins_21,
  input  [63:0] io_ins_22,
  input  [63:0] io_ins_23,
  input  [63:0] io_ins_24,
  input  [63:0] io_ins_25,
  input  [63:0] io_ins_26,
  input  [63:0] io_ins_27,
  input  [63:0] io_ins_28,
  input  [63:0] io_ins_29,
  input  [63:0] io_ins_30,
  input  [63:0] io_ins_31,
  input  [63:0] io_ins_32,
  input  [63:0] io_ins_33,
  input  [63:0] io_ins_34,
  input  [63:0] io_ins_35,
  input  [63:0] io_ins_36,
  input  [63:0] io_ins_37,
  input  [63:0] io_ins_38,
  input  [63:0] io_ins_39,
  input  [63:0] io_ins_40,
  input  [63:0] io_ins_41,
  input  [63:0] io_ins_42,
  input  [63:0] io_ins_43,
  input  [63:0] io_ins_44,
  input  [63:0] io_ins_45,
  input  [63:0] io_ins_46,
  input  [63:0] io_ins_47,
  input  [63:0] io_ins_48,
  input  [63:0] io_ins_49,
  input  [63:0] io_ins_50,
  input  [63:0] io_ins_51,
  input  [63:0] io_ins_52,
  input  [63:0] io_ins_53,
  input  [63:0] io_ins_54,
  input  [63:0] io_ins_55,
  input  [63:0] io_ins_56,
  input  [63:0] io_ins_57,
  input  [63:0] io_ins_58,
  input  [63:0] io_ins_59,
  input  [63:0] io_ins_60,
  input  [63:0] io_ins_61,
  input  [63:0] io_ins_62,
  input  [63:0] io_ins_63,
  input  [63:0] io_ins_64,
  input  [63:0] io_ins_65,
  input  [63:0] io_ins_66,
  input  [63:0] io_ins_67,
  input  [63:0] io_ins_68,
  input  [63:0] io_ins_69,
  input  [63:0] io_ins_70,
  input  [63:0] io_ins_71,
  input  [63:0] io_ins_72,
  input  [63:0] io_ins_73,
  input  [63:0] io_ins_74,
  input  [63:0] io_ins_75,
  input  [63:0] io_ins_76,
  input  [63:0] io_ins_77,
  input  [63:0] io_ins_78,
  input  [63:0] io_ins_79,
  input  [63:0] io_ins_80,
  input  [63:0] io_ins_81,
  input  [63:0] io_ins_82,
  input  [63:0] io_ins_83,
  input  [63:0] io_ins_84,
  input  [63:0] io_ins_85,
  input  [63:0] io_ins_86,
  input  [63:0] io_ins_87,
  input  [63:0] io_ins_88,
  input  [63:0] io_ins_89,
  input  [63:0] io_ins_90,
  input  [63:0] io_ins_91,
  input  [63:0] io_ins_92,
  input  [63:0] io_ins_93,
  input  [63:0] io_ins_94,
  input  [63:0] io_ins_95,
  input  [63:0] io_ins_96,
  input  [63:0] io_ins_97,
  input  [63:0] io_ins_98,
  input  [63:0] io_ins_99,
  input  [63:0] io_ins_100,
  input  [63:0] io_ins_101,
  input  [63:0] io_ins_102,
  input  [63:0] io_ins_103,
  input  [63:0] io_ins_104,
  input  [63:0] io_ins_105,
  input  [63:0] io_ins_106,
  input  [63:0] io_ins_107,
  input  [63:0] io_ins_108,
  input  [63:0] io_ins_109,
  input  [63:0] io_ins_110,
  input  [63:0] io_ins_111,
  input  [63:0] io_ins_112,
  input  [63:0] io_ins_113,
  input  [63:0] io_ins_114,
  input  [63:0] io_ins_115,
  input  [63:0] io_ins_116,
  input  [63:0] io_ins_117,
  input  [63:0] io_ins_118,
  input  [63:0] io_ins_119,
  input  [63:0] io_ins_120,
  input  [63:0] io_ins_121,
  input  [63:0] io_ins_122,
  input  [63:0] io_ins_123,
  input  [63:0] io_ins_124,
  input  [63:0] io_ins_125,
  input  [63:0] io_ins_126,
  input  [63:0] io_ins_127,
  input  [63:0] io_ins_128,
  input  [63:0] io_ins_129,
  input  [63:0] io_ins_130,
  input  [63:0] io_ins_131,
  input  [63:0] io_ins_132,
  input  [63:0] io_ins_133,
  input  [63:0] io_ins_134,
  input  [63:0] io_ins_135,
  input  [63:0] io_ins_136,
  input  [63:0] io_ins_137,
  input  [63:0] io_ins_138,
  input  [63:0] io_ins_139,
  input  [63:0] io_ins_140,
  input  [63:0] io_ins_141,
  input  [63:0] io_ins_142,
  input  [63:0] io_ins_143,
  input  [63:0] io_ins_144,
  input  [63:0] io_ins_145,
  input  [63:0] io_ins_146,
  input  [63:0] io_ins_147,
  input  [63:0] io_ins_148,
  input  [63:0] io_ins_149,
  input  [63:0] io_ins_150,
  input  [63:0] io_ins_151,
  input  [63:0] io_ins_152,
  input  [63:0] io_ins_153,
  input  [63:0] io_ins_154,
  input  [63:0] io_ins_155,
  input  [63:0] io_ins_156,
  input  [63:0] io_ins_157,
  input  [63:0] io_ins_158,
  input  [63:0] io_ins_159,
  input  [63:0] io_ins_160,
  input  [63:0] io_ins_161,
  input  [63:0] io_ins_162,
  input  [63:0] io_ins_163,
  input  [63:0] io_ins_164,
  input  [63:0] io_ins_165,
  input  [63:0] io_ins_166,
  input  [63:0] io_ins_167,
  input  [63:0] io_ins_168,
  input  [63:0] io_ins_169,
  input  [63:0] io_ins_170,
  input  [63:0] io_ins_171,
  input  [63:0] io_ins_172,
  input  [63:0] io_ins_173,
  input  [63:0] io_ins_174,
  input  [63:0] io_ins_175,
  input  [63:0] io_ins_176,
  input  [63:0] io_ins_177,
  input  [63:0] io_ins_178,
  input  [63:0] io_ins_179,
  input  [63:0] io_ins_180,
  input  [63:0] io_ins_181,
  input  [63:0] io_ins_182,
  input  [63:0] io_ins_183,
  input  [63:0] io_ins_184,
  input  [63:0] io_ins_185,
  input  [63:0] io_ins_186,
  input  [63:0] io_ins_187,
  input  [63:0] io_ins_188,
  input  [63:0] io_ins_189,
  input  [63:0] io_ins_190,
  input  [63:0] io_ins_191,
  input  [63:0] io_ins_192,
  input  [63:0] io_ins_193,
  input  [63:0] io_ins_194,
  input  [63:0] io_ins_195,
  input  [63:0] io_ins_196,
  input  [63:0] io_ins_197,
  input  [63:0] io_ins_198,
  input  [63:0] io_ins_199,
  input  [63:0] io_ins_200,
  input  [63:0] io_ins_201,
  input  [63:0] io_ins_202,
  input  [63:0] io_ins_203,
  input  [63:0] io_ins_204,
  input  [63:0] io_ins_205,
  input  [63:0] io_ins_206,
  input  [63:0] io_ins_207,
  input  [63:0] io_ins_208,
  input  [63:0] io_ins_209,
  input  [63:0] io_ins_210,
  input  [63:0] io_ins_211,
  input  [63:0] io_ins_212,
  input  [63:0] io_ins_213,
  input  [63:0] io_ins_214,
  input  [63:0] io_ins_215,
  input  [63:0] io_ins_216,
  input  [63:0] io_ins_217,
  input  [63:0] io_ins_218,
  input  [63:0] io_ins_219,
  input  [63:0] io_ins_220,
  input  [63:0] io_ins_221,
  input  [63:0] io_ins_222,
  input  [63:0] io_ins_223,
  input  [63:0] io_ins_224,
  input  [63:0] io_ins_225,
  input  [63:0] io_ins_226,
  input  [63:0] io_ins_227,
  input  [63:0] io_ins_228,
  input  [63:0] io_ins_229,
  input  [63:0] io_ins_230,
  input  [63:0] io_ins_231,
  input  [63:0] io_ins_232,
  input  [63:0] io_ins_233,
  input  [63:0] io_ins_234,
  input  [63:0] io_ins_235,
  input  [7:0]  io_sel,
  output [63:0] io_out
);
  wire [63:0] _GEN_0;
  wire [63:0] _GEN_1;
  wire [63:0] _GEN_2;
  wire [63:0] _GEN_3;
  wire [63:0] _GEN_4;
  wire [63:0] _GEN_5;
  wire [63:0] _GEN_6;
  wire [63:0] _GEN_7;
  wire [63:0] _GEN_8;
  wire [63:0] _GEN_9;
  wire [63:0] _GEN_10;
  wire [63:0] _GEN_11;
  wire [63:0] _GEN_12;
  wire [63:0] _GEN_13;
  wire [63:0] _GEN_14;
  wire [63:0] _GEN_15;
  wire [63:0] _GEN_16;
  wire [63:0] _GEN_17;
  wire [63:0] _GEN_18;
  wire [63:0] _GEN_19;
  wire [63:0] _GEN_20;
  wire [63:0] _GEN_21;
  wire [63:0] _GEN_22;
  wire [63:0] _GEN_23;
  wire [63:0] _GEN_24;
  wire [63:0] _GEN_25;
  wire [63:0] _GEN_26;
  wire [63:0] _GEN_27;
  wire [63:0] _GEN_28;
  wire [63:0] _GEN_29;
  wire [63:0] _GEN_30;
  wire [63:0] _GEN_31;
  wire [63:0] _GEN_32;
  wire [63:0] _GEN_33;
  wire [63:0] _GEN_34;
  wire [63:0] _GEN_35;
  wire [63:0] _GEN_36;
  wire [63:0] _GEN_37;
  wire [63:0] _GEN_38;
  wire [63:0] _GEN_39;
  wire [63:0] _GEN_40;
  wire [63:0] _GEN_41;
  wire [63:0] _GEN_42;
  wire [63:0] _GEN_43;
  wire [63:0] _GEN_44;
  wire [63:0] _GEN_45;
  wire [63:0] _GEN_46;
  wire [63:0] _GEN_47;
  wire [63:0] _GEN_48;
  wire [63:0] _GEN_49;
  wire [63:0] _GEN_50;
  wire [63:0] _GEN_51;
  wire [63:0] _GEN_52;
  wire [63:0] _GEN_53;
  wire [63:0] _GEN_54;
  wire [63:0] _GEN_55;
  wire [63:0] _GEN_56;
  wire [63:0] _GEN_57;
  wire [63:0] _GEN_58;
  wire [63:0] _GEN_59;
  wire [63:0] _GEN_60;
  wire [63:0] _GEN_61;
  wire [63:0] _GEN_62;
  wire [63:0] _GEN_63;
  wire [63:0] _GEN_64;
  wire [63:0] _GEN_65;
  wire [63:0] _GEN_66;
  wire [63:0] _GEN_67;
  wire [63:0] _GEN_68;
  wire [63:0] _GEN_69;
  wire [63:0] _GEN_70;
  wire [63:0] _GEN_71;
  wire [63:0] _GEN_72;
  wire [63:0] _GEN_73;
  wire [63:0] _GEN_74;
  wire [63:0] _GEN_75;
  wire [63:0] _GEN_76;
  wire [63:0] _GEN_77;
  wire [63:0] _GEN_78;
  wire [63:0] _GEN_79;
  wire [63:0] _GEN_80;
  wire [63:0] _GEN_81;
  wire [63:0] _GEN_82;
  wire [63:0] _GEN_83;
  wire [63:0] _GEN_84;
  wire [63:0] _GEN_85;
  wire [63:0] _GEN_86;
  wire [63:0] _GEN_87;
  wire [63:0] _GEN_88;
  wire [63:0] _GEN_89;
  wire [63:0] _GEN_90;
  wire [63:0] _GEN_91;
  wire [63:0] _GEN_92;
  wire [63:0] _GEN_93;
  wire [63:0] _GEN_94;
  wire [63:0] _GEN_95;
  wire [63:0] _GEN_96;
  wire [63:0] _GEN_97;
  wire [63:0] _GEN_98;
  wire [63:0] _GEN_99;
  wire [63:0] _GEN_100;
  wire [63:0] _GEN_101;
  wire [63:0] _GEN_102;
  wire [63:0] _GEN_103;
  wire [63:0] _GEN_104;
  wire [63:0] _GEN_105;
  wire [63:0] _GEN_106;
  wire [63:0] _GEN_107;
  wire [63:0] _GEN_108;
  wire [63:0] _GEN_109;
  wire [63:0] _GEN_110;
  wire [63:0] _GEN_111;
  wire [63:0] _GEN_112;
  wire [63:0] _GEN_113;
  wire [63:0] _GEN_114;
  wire [63:0] _GEN_115;
  wire [63:0] _GEN_116;
  wire [63:0] _GEN_117;
  wire [63:0] _GEN_118;
  wire [63:0] _GEN_119;
  wire [63:0] _GEN_120;
  wire [63:0] _GEN_121;
  wire [63:0] _GEN_122;
  wire [63:0] _GEN_123;
  wire [63:0] _GEN_124;
  wire [63:0] _GEN_125;
  wire [63:0] _GEN_126;
  wire [63:0] _GEN_127;
  wire [63:0] _GEN_128;
  wire [63:0] _GEN_129;
  wire [63:0] _GEN_130;
  wire [63:0] _GEN_131;
  wire [63:0] _GEN_132;
  wire [63:0] _GEN_133;
  wire [63:0] _GEN_134;
  wire [63:0] _GEN_135;
  wire [63:0] _GEN_136;
  wire [63:0] _GEN_137;
  wire [63:0] _GEN_138;
  wire [63:0] _GEN_139;
  wire [63:0] _GEN_140;
  wire [63:0] _GEN_141;
  wire [63:0] _GEN_142;
  wire [63:0] _GEN_143;
  wire [63:0] _GEN_144;
  wire [63:0] _GEN_145;
  wire [63:0] _GEN_146;
  wire [63:0] _GEN_147;
  wire [63:0] _GEN_148;
  wire [63:0] _GEN_149;
  wire [63:0] _GEN_150;
  wire [63:0] _GEN_151;
  wire [63:0] _GEN_152;
  wire [63:0] _GEN_153;
  wire [63:0] _GEN_154;
  wire [63:0] _GEN_155;
  wire [63:0] _GEN_156;
  wire [63:0] _GEN_157;
  wire [63:0] _GEN_158;
  wire [63:0] _GEN_159;
  wire [63:0] _GEN_160;
  wire [63:0] _GEN_161;
  wire [63:0] _GEN_162;
  wire [63:0] _GEN_163;
  wire [63:0] _GEN_164;
  wire [63:0] _GEN_165;
  wire [63:0] _GEN_166;
  wire [63:0] _GEN_167;
  wire [63:0] _GEN_168;
  wire [63:0] _GEN_169;
  wire [63:0] _GEN_170;
  wire [63:0] _GEN_171;
  wire [63:0] _GEN_172;
  wire [63:0] _GEN_173;
  wire [63:0] _GEN_174;
  wire [63:0] _GEN_175;
  wire [63:0] _GEN_176;
  wire [63:0] _GEN_177;
  wire [63:0] _GEN_178;
  wire [63:0] _GEN_179;
  wire [63:0] _GEN_180;
  wire [63:0] _GEN_181;
  wire [63:0] _GEN_182;
  wire [63:0] _GEN_183;
  wire [63:0] _GEN_184;
  wire [63:0] _GEN_185;
  wire [63:0] _GEN_186;
  wire [63:0] _GEN_187;
  wire [63:0] _GEN_188;
  wire [63:0] _GEN_189;
  wire [63:0] _GEN_190;
  wire [63:0] _GEN_191;
  wire [63:0] _GEN_192;
  wire [63:0] _GEN_193;
  wire [63:0] _GEN_194;
  wire [63:0] _GEN_195;
  wire [63:0] _GEN_196;
  wire [63:0] _GEN_197;
  wire [63:0] _GEN_198;
  wire [63:0] _GEN_199;
  wire [63:0] _GEN_200;
  wire [63:0] _GEN_201;
  wire [63:0] _GEN_202;
  wire [63:0] _GEN_203;
  wire [63:0] _GEN_204;
  wire [63:0] _GEN_205;
  wire [63:0] _GEN_206;
  wire [63:0] _GEN_207;
  wire [63:0] _GEN_208;
  wire [63:0] _GEN_209;
  wire [63:0] _GEN_210;
  wire [63:0] _GEN_211;
  wire [63:0] _GEN_212;
  wire [63:0] _GEN_213;
  wire [63:0] _GEN_214;
  wire [63:0] _GEN_215;
  wire [63:0] _GEN_216;
  wire [63:0] _GEN_217;
  wire [63:0] _GEN_218;
  wire [63:0] _GEN_219;
  wire [63:0] _GEN_220;
  wire [63:0] _GEN_221;
  wire [63:0] _GEN_222;
  wire [63:0] _GEN_223;
  wire [63:0] _GEN_224;
  wire [63:0] _GEN_225;
  wire [63:0] _GEN_226;
  wire [63:0] _GEN_227;
  wire [63:0] _GEN_228;
  wire [63:0] _GEN_229;
  wire [63:0] _GEN_230;
  wire [63:0] _GEN_231;
  wire [63:0] _GEN_232;
  wire [63:0] _GEN_233;
  wire [63:0] _GEN_234;
  wire [63:0] _GEN_235;
  assign _GEN_1 = 8'h1 == io_sel ? io_ins_1 : io_ins_0;
  assign _GEN_2 = 8'h2 == io_sel ? io_ins_2 : _GEN_1;
  assign _GEN_3 = 8'h3 == io_sel ? io_ins_3 : _GEN_2;
  assign _GEN_4 = 8'h4 == io_sel ? io_ins_4 : _GEN_3;
  assign _GEN_5 = 8'h5 == io_sel ? io_ins_5 : _GEN_4;
  assign _GEN_6 = 8'h6 == io_sel ? io_ins_6 : _GEN_5;
  assign _GEN_7 = 8'h7 == io_sel ? io_ins_7 : _GEN_6;
  assign _GEN_8 = 8'h8 == io_sel ? io_ins_8 : _GEN_7;
  assign _GEN_9 = 8'h9 == io_sel ? io_ins_9 : _GEN_8;
  assign _GEN_10 = 8'ha == io_sel ? io_ins_10 : _GEN_9;
  assign _GEN_11 = 8'hb == io_sel ? io_ins_11 : _GEN_10;
  assign _GEN_12 = 8'hc == io_sel ? io_ins_12 : _GEN_11;
  assign _GEN_13 = 8'hd == io_sel ? io_ins_13 : _GEN_12;
  assign _GEN_14 = 8'he == io_sel ? io_ins_14 : _GEN_13;
  assign _GEN_15 = 8'hf == io_sel ? io_ins_15 : _GEN_14;
  assign _GEN_16 = 8'h10 == io_sel ? io_ins_16 : _GEN_15;
  assign _GEN_17 = 8'h11 == io_sel ? io_ins_17 : _GEN_16;
  assign _GEN_18 = 8'h12 == io_sel ? io_ins_18 : _GEN_17;
  assign _GEN_19 = 8'h13 == io_sel ? io_ins_19 : _GEN_18;
  assign _GEN_20 = 8'h14 == io_sel ? io_ins_20 : _GEN_19;
  assign _GEN_21 = 8'h15 == io_sel ? io_ins_21 : _GEN_20;
  assign _GEN_22 = 8'h16 == io_sel ? io_ins_22 : _GEN_21;
  assign _GEN_23 = 8'h17 == io_sel ? io_ins_23 : _GEN_22;
  assign _GEN_24 = 8'h18 == io_sel ? io_ins_24 : _GEN_23;
  assign _GEN_25 = 8'h19 == io_sel ? io_ins_25 : _GEN_24;
  assign _GEN_26 = 8'h1a == io_sel ? io_ins_26 : _GEN_25;
  assign _GEN_27 = 8'h1b == io_sel ? io_ins_27 : _GEN_26;
  assign _GEN_28 = 8'h1c == io_sel ? io_ins_28 : _GEN_27;
  assign _GEN_29 = 8'h1d == io_sel ? io_ins_29 : _GEN_28;
  assign _GEN_30 = 8'h1e == io_sel ? io_ins_30 : _GEN_29;
  assign _GEN_31 = 8'h1f == io_sel ? io_ins_31 : _GEN_30;
  assign _GEN_32 = 8'h20 == io_sel ? io_ins_32 : _GEN_31;
  assign _GEN_33 = 8'h21 == io_sel ? io_ins_33 : _GEN_32;
  assign _GEN_34 = 8'h22 == io_sel ? io_ins_34 : _GEN_33;
  assign _GEN_35 = 8'h23 == io_sel ? io_ins_35 : _GEN_34;
  assign _GEN_36 = 8'h24 == io_sel ? io_ins_36 : _GEN_35;
  assign _GEN_37 = 8'h25 == io_sel ? io_ins_37 : _GEN_36;
  assign _GEN_38 = 8'h26 == io_sel ? io_ins_38 : _GEN_37;
  assign _GEN_39 = 8'h27 == io_sel ? io_ins_39 : _GEN_38;
  assign _GEN_40 = 8'h28 == io_sel ? io_ins_40 : _GEN_39;
  assign _GEN_41 = 8'h29 == io_sel ? io_ins_41 : _GEN_40;
  assign _GEN_42 = 8'h2a == io_sel ? io_ins_42 : _GEN_41;
  assign _GEN_43 = 8'h2b == io_sel ? io_ins_43 : _GEN_42;
  assign _GEN_44 = 8'h2c == io_sel ? io_ins_44 : _GEN_43;
  assign _GEN_45 = 8'h2d == io_sel ? io_ins_45 : _GEN_44;
  assign _GEN_46 = 8'h2e == io_sel ? io_ins_46 : _GEN_45;
  assign _GEN_47 = 8'h2f == io_sel ? io_ins_47 : _GEN_46;
  assign _GEN_48 = 8'h30 == io_sel ? io_ins_48 : _GEN_47;
  assign _GEN_49 = 8'h31 == io_sel ? io_ins_49 : _GEN_48;
  assign _GEN_50 = 8'h32 == io_sel ? io_ins_50 : _GEN_49;
  assign _GEN_51 = 8'h33 == io_sel ? io_ins_51 : _GEN_50;
  assign _GEN_52 = 8'h34 == io_sel ? io_ins_52 : _GEN_51;
  assign _GEN_53 = 8'h35 == io_sel ? io_ins_53 : _GEN_52;
  assign _GEN_54 = 8'h36 == io_sel ? io_ins_54 : _GEN_53;
  assign _GEN_55 = 8'h37 == io_sel ? io_ins_55 : _GEN_54;
  assign _GEN_56 = 8'h38 == io_sel ? io_ins_56 : _GEN_55;
  assign _GEN_57 = 8'h39 == io_sel ? io_ins_57 : _GEN_56;
  assign _GEN_58 = 8'h3a == io_sel ? io_ins_58 : _GEN_57;
  assign _GEN_59 = 8'h3b == io_sel ? io_ins_59 : _GEN_58;
  assign _GEN_60 = 8'h3c == io_sel ? io_ins_60 : _GEN_59;
  assign _GEN_61 = 8'h3d == io_sel ? io_ins_61 : _GEN_60;
  assign _GEN_62 = 8'h3e == io_sel ? io_ins_62 : _GEN_61;
  assign _GEN_63 = 8'h3f == io_sel ? io_ins_63 : _GEN_62;
  assign _GEN_64 = 8'h40 == io_sel ? io_ins_64 : _GEN_63;
  assign _GEN_65 = 8'h41 == io_sel ? io_ins_65 : _GEN_64;
  assign _GEN_66 = 8'h42 == io_sel ? io_ins_66 : _GEN_65;
  assign _GEN_67 = 8'h43 == io_sel ? io_ins_67 : _GEN_66;
  assign _GEN_68 = 8'h44 == io_sel ? io_ins_68 : _GEN_67;
  assign _GEN_69 = 8'h45 == io_sel ? io_ins_69 : _GEN_68;
  assign _GEN_70 = 8'h46 == io_sel ? io_ins_70 : _GEN_69;
  assign _GEN_71 = 8'h47 == io_sel ? io_ins_71 : _GEN_70;
  assign _GEN_72 = 8'h48 == io_sel ? io_ins_72 : _GEN_71;
  assign _GEN_73 = 8'h49 == io_sel ? io_ins_73 : _GEN_72;
  assign _GEN_74 = 8'h4a == io_sel ? io_ins_74 : _GEN_73;
  assign _GEN_75 = 8'h4b == io_sel ? io_ins_75 : _GEN_74;
  assign _GEN_76 = 8'h4c == io_sel ? io_ins_76 : _GEN_75;
  assign _GEN_77 = 8'h4d == io_sel ? io_ins_77 : _GEN_76;
  assign _GEN_78 = 8'h4e == io_sel ? io_ins_78 : _GEN_77;
  assign _GEN_79 = 8'h4f == io_sel ? io_ins_79 : _GEN_78;
  assign _GEN_80 = 8'h50 == io_sel ? io_ins_80 : _GEN_79;
  assign _GEN_81 = 8'h51 == io_sel ? io_ins_81 : _GEN_80;
  assign _GEN_82 = 8'h52 == io_sel ? io_ins_82 : _GEN_81;
  assign _GEN_83 = 8'h53 == io_sel ? io_ins_83 : _GEN_82;
  assign _GEN_84 = 8'h54 == io_sel ? io_ins_84 : _GEN_83;
  assign _GEN_85 = 8'h55 == io_sel ? io_ins_85 : _GEN_84;
  assign _GEN_86 = 8'h56 == io_sel ? io_ins_86 : _GEN_85;
  assign _GEN_87 = 8'h57 == io_sel ? io_ins_87 : _GEN_86;
  assign _GEN_88 = 8'h58 == io_sel ? io_ins_88 : _GEN_87;
  assign _GEN_89 = 8'h59 == io_sel ? io_ins_89 : _GEN_88;
  assign _GEN_90 = 8'h5a == io_sel ? io_ins_90 : _GEN_89;
  assign _GEN_91 = 8'h5b == io_sel ? io_ins_91 : _GEN_90;
  assign _GEN_92 = 8'h5c == io_sel ? io_ins_92 : _GEN_91;
  assign _GEN_93 = 8'h5d == io_sel ? io_ins_93 : _GEN_92;
  assign _GEN_94 = 8'h5e == io_sel ? io_ins_94 : _GEN_93;
  assign _GEN_95 = 8'h5f == io_sel ? io_ins_95 : _GEN_94;
  assign _GEN_96 = 8'h60 == io_sel ? io_ins_96 : _GEN_95;
  assign _GEN_97 = 8'h61 == io_sel ? io_ins_97 : _GEN_96;
  assign _GEN_98 = 8'h62 == io_sel ? io_ins_98 : _GEN_97;
  assign _GEN_99 = 8'h63 == io_sel ? io_ins_99 : _GEN_98;
  assign _GEN_100 = 8'h64 == io_sel ? io_ins_100 : _GEN_99;
  assign _GEN_101 = 8'h65 == io_sel ? io_ins_101 : _GEN_100;
  assign _GEN_102 = 8'h66 == io_sel ? io_ins_102 : _GEN_101;
  assign _GEN_103 = 8'h67 == io_sel ? io_ins_103 : _GEN_102;
  assign _GEN_104 = 8'h68 == io_sel ? io_ins_104 : _GEN_103;
  assign _GEN_105 = 8'h69 == io_sel ? io_ins_105 : _GEN_104;
  assign _GEN_106 = 8'h6a == io_sel ? io_ins_106 : _GEN_105;
  assign _GEN_107 = 8'h6b == io_sel ? io_ins_107 : _GEN_106;
  assign _GEN_108 = 8'h6c == io_sel ? io_ins_108 : _GEN_107;
  assign _GEN_109 = 8'h6d == io_sel ? io_ins_109 : _GEN_108;
  assign _GEN_110 = 8'h6e == io_sel ? io_ins_110 : _GEN_109;
  assign _GEN_111 = 8'h6f == io_sel ? io_ins_111 : _GEN_110;
  assign _GEN_112 = 8'h70 == io_sel ? io_ins_112 : _GEN_111;
  assign _GEN_113 = 8'h71 == io_sel ? io_ins_113 : _GEN_112;
  assign _GEN_114 = 8'h72 == io_sel ? io_ins_114 : _GEN_113;
  assign _GEN_115 = 8'h73 == io_sel ? io_ins_115 : _GEN_114;
  assign _GEN_116 = 8'h74 == io_sel ? io_ins_116 : _GEN_115;
  assign _GEN_117 = 8'h75 == io_sel ? io_ins_117 : _GEN_116;
  assign _GEN_118 = 8'h76 == io_sel ? io_ins_118 : _GEN_117;
  assign _GEN_119 = 8'h77 == io_sel ? io_ins_119 : _GEN_118;
  assign _GEN_120 = 8'h78 == io_sel ? io_ins_120 : _GEN_119;
  assign _GEN_121 = 8'h79 == io_sel ? io_ins_121 : _GEN_120;
  assign _GEN_122 = 8'h7a == io_sel ? io_ins_122 : _GEN_121;
  assign _GEN_123 = 8'h7b == io_sel ? io_ins_123 : _GEN_122;
  assign _GEN_124 = 8'h7c == io_sel ? io_ins_124 : _GEN_123;
  assign _GEN_125 = 8'h7d == io_sel ? io_ins_125 : _GEN_124;
  assign _GEN_126 = 8'h7e == io_sel ? io_ins_126 : _GEN_125;
  assign _GEN_127 = 8'h7f == io_sel ? io_ins_127 : _GEN_126;
  assign _GEN_128 = 8'h80 == io_sel ? io_ins_128 : _GEN_127;
  assign _GEN_129 = 8'h81 == io_sel ? io_ins_129 : _GEN_128;
  assign _GEN_130 = 8'h82 == io_sel ? io_ins_130 : _GEN_129;
  assign _GEN_131 = 8'h83 == io_sel ? io_ins_131 : _GEN_130;
  assign _GEN_132 = 8'h84 == io_sel ? io_ins_132 : _GEN_131;
  assign _GEN_133 = 8'h85 == io_sel ? io_ins_133 : _GEN_132;
  assign _GEN_134 = 8'h86 == io_sel ? io_ins_134 : _GEN_133;
  assign _GEN_135 = 8'h87 == io_sel ? io_ins_135 : _GEN_134;
  assign _GEN_136 = 8'h88 == io_sel ? io_ins_136 : _GEN_135;
  assign _GEN_137 = 8'h89 == io_sel ? io_ins_137 : _GEN_136;
  assign _GEN_138 = 8'h8a == io_sel ? io_ins_138 : _GEN_137;
  assign _GEN_139 = 8'h8b == io_sel ? io_ins_139 : _GEN_138;
  assign _GEN_140 = 8'h8c == io_sel ? io_ins_140 : _GEN_139;
  assign _GEN_141 = 8'h8d == io_sel ? io_ins_141 : _GEN_140;
  assign _GEN_142 = 8'h8e == io_sel ? io_ins_142 : _GEN_141;
  assign _GEN_143 = 8'h8f == io_sel ? io_ins_143 : _GEN_142;
  assign _GEN_144 = 8'h90 == io_sel ? io_ins_144 : _GEN_143;
  assign _GEN_145 = 8'h91 == io_sel ? io_ins_145 : _GEN_144;
  assign _GEN_146 = 8'h92 == io_sel ? io_ins_146 : _GEN_145;
  assign _GEN_147 = 8'h93 == io_sel ? io_ins_147 : _GEN_146;
  assign _GEN_148 = 8'h94 == io_sel ? io_ins_148 : _GEN_147;
  assign _GEN_149 = 8'h95 == io_sel ? io_ins_149 : _GEN_148;
  assign _GEN_150 = 8'h96 == io_sel ? io_ins_150 : _GEN_149;
  assign _GEN_151 = 8'h97 == io_sel ? io_ins_151 : _GEN_150;
  assign _GEN_152 = 8'h98 == io_sel ? io_ins_152 : _GEN_151;
  assign _GEN_153 = 8'h99 == io_sel ? io_ins_153 : _GEN_152;
  assign _GEN_154 = 8'h9a == io_sel ? io_ins_154 : _GEN_153;
  assign _GEN_155 = 8'h9b == io_sel ? io_ins_155 : _GEN_154;
  assign _GEN_156 = 8'h9c == io_sel ? io_ins_156 : _GEN_155;
  assign _GEN_157 = 8'h9d == io_sel ? io_ins_157 : _GEN_156;
  assign _GEN_158 = 8'h9e == io_sel ? io_ins_158 : _GEN_157;
  assign _GEN_159 = 8'h9f == io_sel ? io_ins_159 : _GEN_158;
  assign _GEN_160 = 8'ha0 == io_sel ? io_ins_160 : _GEN_159;
  assign _GEN_161 = 8'ha1 == io_sel ? io_ins_161 : _GEN_160;
  assign _GEN_162 = 8'ha2 == io_sel ? io_ins_162 : _GEN_161;
  assign _GEN_163 = 8'ha3 == io_sel ? io_ins_163 : _GEN_162;
  assign _GEN_164 = 8'ha4 == io_sel ? io_ins_164 : _GEN_163;
  assign _GEN_165 = 8'ha5 == io_sel ? io_ins_165 : _GEN_164;
  assign _GEN_166 = 8'ha6 == io_sel ? io_ins_166 : _GEN_165;
  assign _GEN_167 = 8'ha7 == io_sel ? io_ins_167 : _GEN_166;
  assign _GEN_168 = 8'ha8 == io_sel ? io_ins_168 : _GEN_167;
  assign _GEN_169 = 8'ha9 == io_sel ? io_ins_169 : _GEN_168;
  assign _GEN_170 = 8'haa == io_sel ? io_ins_170 : _GEN_169;
  assign _GEN_171 = 8'hab == io_sel ? io_ins_171 : _GEN_170;
  assign _GEN_172 = 8'hac == io_sel ? io_ins_172 : _GEN_171;
  assign _GEN_173 = 8'had == io_sel ? io_ins_173 : _GEN_172;
  assign _GEN_174 = 8'hae == io_sel ? io_ins_174 : _GEN_173;
  assign _GEN_175 = 8'haf == io_sel ? io_ins_175 : _GEN_174;
  assign _GEN_176 = 8'hb0 == io_sel ? io_ins_176 : _GEN_175;
  assign _GEN_177 = 8'hb1 == io_sel ? io_ins_177 : _GEN_176;
  assign _GEN_178 = 8'hb2 == io_sel ? io_ins_178 : _GEN_177;
  assign _GEN_179 = 8'hb3 == io_sel ? io_ins_179 : _GEN_178;
  assign _GEN_180 = 8'hb4 == io_sel ? io_ins_180 : _GEN_179;
  assign _GEN_181 = 8'hb5 == io_sel ? io_ins_181 : _GEN_180;
  assign _GEN_182 = 8'hb6 == io_sel ? io_ins_182 : _GEN_181;
  assign _GEN_183 = 8'hb7 == io_sel ? io_ins_183 : _GEN_182;
  assign _GEN_184 = 8'hb8 == io_sel ? io_ins_184 : _GEN_183;
  assign _GEN_185 = 8'hb9 == io_sel ? io_ins_185 : _GEN_184;
  assign _GEN_186 = 8'hba == io_sel ? io_ins_186 : _GEN_185;
  assign _GEN_187 = 8'hbb == io_sel ? io_ins_187 : _GEN_186;
  assign _GEN_188 = 8'hbc == io_sel ? io_ins_188 : _GEN_187;
  assign _GEN_189 = 8'hbd == io_sel ? io_ins_189 : _GEN_188;
  assign _GEN_190 = 8'hbe == io_sel ? io_ins_190 : _GEN_189;
  assign _GEN_191 = 8'hbf == io_sel ? io_ins_191 : _GEN_190;
  assign _GEN_192 = 8'hc0 == io_sel ? io_ins_192 : _GEN_191;
  assign _GEN_193 = 8'hc1 == io_sel ? io_ins_193 : _GEN_192;
  assign _GEN_194 = 8'hc2 == io_sel ? io_ins_194 : _GEN_193;
  assign _GEN_195 = 8'hc3 == io_sel ? io_ins_195 : _GEN_194;
  assign _GEN_196 = 8'hc4 == io_sel ? io_ins_196 : _GEN_195;
  assign _GEN_197 = 8'hc5 == io_sel ? io_ins_197 : _GEN_196;
  assign _GEN_198 = 8'hc6 == io_sel ? io_ins_198 : _GEN_197;
  assign _GEN_199 = 8'hc7 == io_sel ? io_ins_199 : _GEN_198;
  assign _GEN_200 = 8'hc8 == io_sel ? io_ins_200 : _GEN_199;
  assign _GEN_201 = 8'hc9 == io_sel ? io_ins_201 : _GEN_200;
  assign _GEN_202 = 8'hca == io_sel ? io_ins_202 : _GEN_201;
  assign _GEN_203 = 8'hcb == io_sel ? io_ins_203 : _GEN_202;
  assign _GEN_204 = 8'hcc == io_sel ? io_ins_204 : _GEN_203;
  assign _GEN_205 = 8'hcd == io_sel ? io_ins_205 : _GEN_204;
  assign _GEN_206 = 8'hce == io_sel ? io_ins_206 : _GEN_205;
  assign _GEN_207 = 8'hcf == io_sel ? io_ins_207 : _GEN_206;
  assign _GEN_208 = 8'hd0 == io_sel ? io_ins_208 : _GEN_207;
  assign _GEN_209 = 8'hd1 == io_sel ? io_ins_209 : _GEN_208;
  assign _GEN_210 = 8'hd2 == io_sel ? io_ins_210 : _GEN_209;
  assign _GEN_211 = 8'hd3 == io_sel ? io_ins_211 : _GEN_210;
  assign _GEN_212 = 8'hd4 == io_sel ? io_ins_212 : _GEN_211;
  assign _GEN_213 = 8'hd5 == io_sel ? io_ins_213 : _GEN_212;
  assign _GEN_214 = 8'hd6 == io_sel ? io_ins_214 : _GEN_213;
  assign _GEN_215 = 8'hd7 == io_sel ? io_ins_215 : _GEN_214;
  assign _GEN_216 = 8'hd8 == io_sel ? io_ins_216 : _GEN_215;
  assign _GEN_217 = 8'hd9 == io_sel ? io_ins_217 : _GEN_216;
  assign _GEN_218 = 8'hda == io_sel ? io_ins_218 : _GEN_217;
  assign _GEN_219 = 8'hdb == io_sel ? io_ins_219 : _GEN_218;
  assign _GEN_220 = 8'hdc == io_sel ? io_ins_220 : _GEN_219;
  assign _GEN_221 = 8'hdd == io_sel ? io_ins_221 : _GEN_220;
  assign _GEN_222 = 8'hde == io_sel ? io_ins_222 : _GEN_221;
  assign _GEN_223 = 8'hdf == io_sel ? io_ins_223 : _GEN_222;
  assign _GEN_224 = 8'he0 == io_sel ? io_ins_224 : _GEN_223;
  assign _GEN_225 = 8'he1 == io_sel ? io_ins_225 : _GEN_224;
  assign _GEN_226 = 8'he2 == io_sel ? io_ins_226 : _GEN_225;
  assign _GEN_227 = 8'he3 == io_sel ? io_ins_227 : _GEN_226;
  assign _GEN_228 = 8'he4 == io_sel ? io_ins_228 : _GEN_227;
  assign _GEN_229 = 8'he5 == io_sel ? io_ins_229 : _GEN_228;
  assign _GEN_230 = 8'he6 == io_sel ? io_ins_230 : _GEN_229;
  assign _GEN_231 = 8'he7 == io_sel ? io_ins_231 : _GEN_230;
  assign _GEN_232 = 8'he8 == io_sel ? io_ins_232 : _GEN_231;
  assign _GEN_233 = 8'he9 == io_sel ? io_ins_233 : _GEN_232;
  assign _GEN_234 = 8'hea == io_sel ? io_ins_234 : _GEN_233;
  assign _GEN_235 = 8'heb == io_sel ? io_ins_235 : _GEN_234;
  assign io_out = _GEN_0;
  assign _GEN_0 = _GEN_235;
endmodule
module RegFile(
  input         clock,
  input         reset,
  input  [7:0]  io_raddr,
  input         io_wen,
  input  [7:0]  io_waddr,
  input  [63:0] io_wdata,
  output [63:0] io_rdata,
  output [63:0] io_argIns_0,
  output [63:0] io_argIns_1,
  output [63:0] io_argIns_2,
  input         io_argOuts_0_valid,
  input  [63:0] io_argOuts_0_bits,
  input         io_argOuts_1_valid,
  input  [63:0] io_argOuts_1_bits,
  input  [63:0] io_argOuts_2_bits,
  input  [63:0] io_argOuts_3_bits,
  input  [63:0] io_argOuts_4_bits,
  input  [63:0] io_argOuts_5_bits,
  input  [63:0] io_argOuts_6_bits,
  input  [63:0] io_argOuts_7_bits,
  input  [63:0] io_argOuts_8_bits,
  input  [63:0] io_argOuts_9_bits,
  input  [63:0] io_argOuts_10_bits,
  input  [63:0] io_argOuts_11_bits,
  input  [63:0] io_argOuts_12_bits,
  input  [63:0] io_argOuts_13_bits,
  input  [63:0] io_argOuts_14_bits,
  input  [63:0] io_argOuts_15_bits,
  input  [63:0] io_argOuts_16_bits,
  input  [63:0] io_argOuts_17_bits,
  input  [63:0] io_argOuts_18_bits,
  input  [63:0] io_argOuts_19_bits,
  input  [63:0] io_argOuts_20_bits,
  input  [63:0] io_argOuts_21_bits,
  input  [63:0] io_argOuts_22_bits,
  input  [63:0] io_argOuts_23_bits,
  input  [63:0] io_argOuts_24_bits,
  input  [63:0] io_argOuts_25_bits,
  input  [63:0] io_argOuts_26_bits,
  input  [63:0] io_argOuts_27_bits,
  input  [63:0] io_argOuts_28_bits,
  input  [63:0] io_argOuts_29_bits,
  input  [63:0] io_argOuts_30_bits,
  input  [63:0] io_argOuts_31_bits,
  input  [63:0] io_argOuts_32_bits,
  input  [63:0] io_argOuts_33_bits,
  input  [63:0] io_argOuts_34_bits,
  input  [63:0] io_argOuts_35_bits,
  input  [63:0] io_argOuts_36_bits,
  input  [63:0] io_argOuts_37_bits,
  input  [63:0] io_argOuts_38_bits,
  input  [63:0] io_argOuts_39_bits,
  input  [63:0] io_argOuts_40_bits,
  input  [63:0] io_argOuts_41_bits,
  input  [63:0] io_argOuts_42_bits,
  input  [63:0] io_argOuts_43_bits,
  input  [63:0] io_argOuts_44_bits,
  input  [63:0] io_argOuts_45_bits,
  input  [63:0] io_argOuts_46_bits,
  input  [63:0] io_argOuts_47_bits,
  input  [63:0] io_argOuts_48_bits,
  input  [63:0] io_argOuts_49_bits,
  input  [63:0] io_argOuts_50_bits,
  input  [63:0] io_argOuts_51_bits,
  input  [63:0] io_argOuts_52_bits,
  input  [63:0] io_argOuts_53_bits,
  input  [63:0] io_argOuts_54_bits,
  input  [63:0] io_argOuts_55_bits,
  input  [63:0] io_argOuts_56_bits,
  input  [63:0] io_argOuts_57_bits,
  input  [63:0] io_argOuts_58_bits,
  input  [63:0] io_argOuts_59_bits,
  input  [63:0] io_argOuts_60_bits
);
  wire  regs_0_clock;
  wire  regs_0_reset;
  wire [63:0] regs_0_io_in;
  wire [63:0] regs_0_io_init;
  wire [63:0] regs_0_io_out;
  wire  regs_0_io_enable;
  wire  _T_731;
  wire  _T_732;
  wire  regs_1_clock;
  wire  regs_1_reset;
  wire [63:0] regs_1_io_in;
  wire [63:0] regs_1_io_init;
  wire [63:0] regs_1_io_out;
  wire  regs_1_io_enable;
  wire  _T_735;
  wire  _T_736;
  wire  _T_740;
  wire [63:0] _T_744;
  wire  regs_2_clock;
  wire  regs_2_reset;
  wire [63:0] regs_2_io_in;
  wire [63:0] regs_2_io_init;
  wire [63:0] regs_2_io_out;
  wire  regs_2_io_enable;
  wire  _T_747;
  wire  _T_748;
  wire  regs_3_clock;
  wire  regs_3_reset;
  wire [63:0] regs_3_io_in;
  wire [63:0] regs_3_io_init;
  wire [63:0] regs_3_io_out;
  wire  regs_3_io_enable;
  wire  _T_751;
  wire  _T_752;
  wire  _T_753;
  wire [63:0] _T_754;
  wire  regs_4_clock;
  wire  regs_4_reset;
  wire [63:0] regs_4_io_in;
  wire [63:0] regs_4_io_init;
  wire [63:0] regs_4_io_out;
  wire  regs_4_io_enable;
  wire  regs_5_clock;
  wire  regs_5_reset;
  wire [63:0] regs_5_io_in;
  wire [63:0] regs_5_io_init;
  wire [63:0] regs_5_io_out;
  wire  regs_5_io_enable;
  wire  regs_6_clock;
  wire  regs_6_reset;
  wire [63:0] regs_6_io_in;
  wire [63:0] regs_6_io_init;
  wire [63:0] regs_6_io_out;
  wire  regs_6_io_enable;
  wire  regs_7_clock;
  wire  regs_7_reset;
  wire [63:0] regs_7_io_in;
  wire [63:0] regs_7_io_init;
  wire [63:0] regs_7_io_out;
  wire  regs_7_io_enable;
  wire  regs_8_clock;
  wire  regs_8_reset;
  wire [63:0] regs_8_io_in;
  wire [63:0] regs_8_io_init;
  wire [63:0] regs_8_io_out;
  wire  regs_8_io_enable;
  wire  regs_9_clock;
  wire  regs_9_reset;
  wire [63:0] regs_9_io_in;
  wire [63:0] regs_9_io_init;
  wire [63:0] regs_9_io_out;
  wire  regs_9_io_enable;
  wire  regs_10_clock;
  wire  regs_10_reset;
  wire [63:0] regs_10_io_in;
  wire [63:0] regs_10_io_init;
  wire [63:0] regs_10_io_out;
  wire  regs_10_io_enable;
  wire  regs_11_clock;
  wire  regs_11_reset;
  wire [63:0] regs_11_io_in;
  wire [63:0] regs_11_io_init;
  wire [63:0] regs_11_io_out;
  wire  regs_11_io_enable;
  wire  regs_12_clock;
  wire  regs_12_reset;
  wire [63:0] regs_12_io_in;
  wire [63:0] regs_12_io_init;
  wire [63:0] regs_12_io_out;
  wire  regs_12_io_enable;
  wire  regs_13_clock;
  wire  regs_13_reset;
  wire [63:0] regs_13_io_in;
  wire [63:0] regs_13_io_init;
  wire [63:0] regs_13_io_out;
  wire  regs_13_io_enable;
  wire  regs_14_clock;
  wire  regs_14_reset;
  wire [63:0] regs_14_io_in;
  wire [63:0] regs_14_io_init;
  wire [63:0] regs_14_io_out;
  wire  regs_14_io_enable;
  wire  regs_15_clock;
  wire  regs_15_reset;
  wire [63:0] regs_15_io_in;
  wire [63:0] regs_15_io_init;
  wire [63:0] regs_15_io_out;
  wire  regs_15_io_enable;
  wire  regs_16_clock;
  wire  regs_16_reset;
  wire [63:0] regs_16_io_in;
  wire [63:0] regs_16_io_init;
  wire [63:0] regs_16_io_out;
  wire  regs_16_io_enable;
  wire  regs_17_clock;
  wire  regs_17_reset;
  wire [63:0] regs_17_io_in;
  wire [63:0] regs_17_io_init;
  wire [63:0] regs_17_io_out;
  wire  regs_17_io_enable;
  wire  regs_18_clock;
  wire  regs_18_reset;
  wire [63:0] regs_18_io_in;
  wire [63:0] regs_18_io_init;
  wire [63:0] regs_18_io_out;
  wire  regs_18_io_enable;
  wire  regs_19_clock;
  wire  regs_19_reset;
  wire [63:0] regs_19_io_in;
  wire [63:0] regs_19_io_init;
  wire [63:0] regs_19_io_out;
  wire  regs_19_io_enable;
  wire  regs_20_clock;
  wire  regs_20_reset;
  wire [63:0] regs_20_io_in;
  wire [63:0] regs_20_io_init;
  wire [63:0] regs_20_io_out;
  wire  regs_20_io_enable;
  wire  regs_21_clock;
  wire  regs_21_reset;
  wire [63:0] regs_21_io_in;
  wire [63:0] regs_21_io_init;
  wire [63:0] regs_21_io_out;
  wire  regs_21_io_enable;
  wire  regs_22_clock;
  wire  regs_22_reset;
  wire [63:0] regs_22_io_in;
  wire [63:0] regs_22_io_init;
  wire [63:0] regs_22_io_out;
  wire  regs_22_io_enable;
  wire  regs_23_clock;
  wire  regs_23_reset;
  wire [63:0] regs_23_io_in;
  wire [63:0] regs_23_io_init;
  wire [63:0] regs_23_io_out;
  wire  regs_23_io_enable;
  wire  regs_24_clock;
  wire  regs_24_reset;
  wire [63:0] regs_24_io_in;
  wire [63:0] regs_24_io_init;
  wire [63:0] regs_24_io_out;
  wire  regs_24_io_enable;
  wire  regs_25_clock;
  wire  regs_25_reset;
  wire [63:0] regs_25_io_in;
  wire [63:0] regs_25_io_init;
  wire [63:0] regs_25_io_out;
  wire  regs_25_io_enable;
  wire  regs_26_clock;
  wire  regs_26_reset;
  wire [63:0] regs_26_io_in;
  wire [63:0] regs_26_io_init;
  wire [63:0] regs_26_io_out;
  wire  regs_26_io_enable;
  wire  regs_27_clock;
  wire  regs_27_reset;
  wire [63:0] regs_27_io_in;
  wire [63:0] regs_27_io_init;
  wire [63:0] regs_27_io_out;
  wire  regs_27_io_enable;
  wire  regs_28_clock;
  wire  regs_28_reset;
  wire [63:0] regs_28_io_in;
  wire [63:0] regs_28_io_init;
  wire [63:0] regs_28_io_out;
  wire  regs_28_io_enable;
  wire  regs_29_clock;
  wire  regs_29_reset;
  wire [63:0] regs_29_io_in;
  wire [63:0] regs_29_io_init;
  wire [63:0] regs_29_io_out;
  wire  regs_29_io_enable;
  wire  regs_30_clock;
  wire  regs_30_reset;
  wire [63:0] regs_30_io_in;
  wire [63:0] regs_30_io_init;
  wire [63:0] regs_30_io_out;
  wire  regs_30_io_enable;
  wire  regs_31_clock;
  wire  regs_31_reset;
  wire [63:0] regs_31_io_in;
  wire [63:0] regs_31_io_init;
  wire [63:0] regs_31_io_out;
  wire  regs_31_io_enable;
  wire  regs_32_clock;
  wire  regs_32_reset;
  wire [63:0] regs_32_io_in;
  wire [63:0] regs_32_io_init;
  wire [63:0] regs_32_io_out;
  wire  regs_32_io_enable;
  wire  regs_33_clock;
  wire  regs_33_reset;
  wire [63:0] regs_33_io_in;
  wire [63:0] regs_33_io_init;
  wire [63:0] regs_33_io_out;
  wire  regs_33_io_enable;
  wire  regs_34_clock;
  wire  regs_34_reset;
  wire [63:0] regs_34_io_in;
  wire [63:0] regs_34_io_init;
  wire [63:0] regs_34_io_out;
  wire  regs_34_io_enable;
  wire  regs_35_clock;
  wire  regs_35_reset;
  wire [63:0] regs_35_io_in;
  wire [63:0] regs_35_io_init;
  wire [63:0] regs_35_io_out;
  wire  regs_35_io_enable;
  wire  regs_36_clock;
  wire  regs_36_reset;
  wire [63:0] regs_36_io_in;
  wire [63:0] regs_36_io_init;
  wire [63:0] regs_36_io_out;
  wire  regs_36_io_enable;
  wire  regs_37_clock;
  wire  regs_37_reset;
  wire [63:0] regs_37_io_in;
  wire [63:0] regs_37_io_init;
  wire [63:0] regs_37_io_out;
  wire  regs_37_io_enable;
  wire  regs_38_clock;
  wire  regs_38_reset;
  wire [63:0] regs_38_io_in;
  wire [63:0] regs_38_io_init;
  wire [63:0] regs_38_io_out;
  wire  regs_38_io_enable;
  wire  regs_39_clock;
  wire  regs_39_reset;
  wire [63:0] regs_39_io_in;
  wire [63:0] regs_39_io_init;
  wire [63:0] regs_39_io_out;
  wire  regs_39_io_enable;
  wire  regs_40_clock;
  wire  regs_40_reset;
  wire [63:0] regs_40_io_in;
  wire [63:0] regs_40_io_init;
  wire [63:0] regs_40_io_out;
  wire  regs_40_io_enable;
  wire  regs_41_clock;
  wire  regs_41_reset;
  wire [63:0] regs_41_io_in;
  wire [63:0] regs_41_io_init;
  wire [63:0] regs_41_io_out;
  wire  regs_41_io_enable;
  wire  regs_42_clock;
  wire  regs_42_reset;
  wire [63:0] regs_42_io_in;
  wire [63:0] regs_42_io_init;
  wire [63:0] regs_42_io_out;
  wire  regs_42_io_enable;
  wire  regs_43_clock;
  wire  regs_43_reset;
  wire [63:0] regs_43_io_in;
  wire [63:0] regs_43_io_init;
  wire [63:0] regs_43_io_out;
  wire  regs_43_io_enable;
  wire  regs_44_clock;
  wire  regs_44_reset;
  wire [63:0] regs_44_io_in;
  wire [63:0] regs_44_io_init;
  wire [63:0] regs_44_io_out;
  wire  regs_44_io_enable;
  wire  regs_45_clock;
  wire  regs_45_reset;
  wire [63:0] regs_45_io_in;
  wire [63:0] regs_45_io_init;
  wire [63:0] regs_45_io_out;
  wire  regs_45_io_enable;
  wire  regs_46_clock;
  wire  regs_46_reset;
  wire [63:0] regs_46_io_in;
  wire [63:0] regs_46_io_init;
  wire [63:0] regs_46_io_out;
  wire  regs_46_io_enable;
  wire  regs_47_clock;
  wire  regs_47_reset;
  wire [63:0] regs_47_io_in;
  wire [63:0] regs_47_io_init;
  wire [63:0] regs_47_io_out;
  wire  regs_47_io_enable;
  wire  regs_48_clock;
  wire  regs_48_reset;
  wire [63:0] regs_48_io_in;
  wire [63:0] regs_48_io_init;
  wire [63:0] regs_48_io_out;
  wire  regs_48_io_enable;
  wire  regs_49_clock;
  wire  regs_49_reset;
  wire [63:0] regs_49_io_in;
  wire [63:0] regs_49_io_init;
  wire [63:0] regs_49_io_out;
  wire  regs_49_io_enable;
  wire  regs_50_clock;
  wire  regs_50_reset;
  wire [63:0] regs_50_io_in;
  wire [63:0] regs_50_io_init;
  wire [63:0] regs_50_io_out;
  wire  regs_50_io_enable;
  wire  regs_51_clock;
  wire  regs_51_reset;
  wire [63:0] regs_51_io_in;
  wire [63:0] regs_51_io_init;
  wire [63:0] regs_51_io_out;
  wire  regs_51_io_enable;
  wire  regs_52_clock;
  wire  regs_52_reset;
  wire [63:0] regs_52_io_in;
  wire [63:0] regs_52_io_init;
  wire [63:0] regs_52_io_out;
  wire  regs_52_io_enable;
  wire  regs_53_clock;
  wire  regs_53_reset;
  wire [63:0] regs_53_io_in;
  wire [63:0] regs_53_io_init;
  wire [63:0] regs_53_io_out;
  wire  regs_53_io_enable;
  wire  regs_54_clock;
  wire  regs_54_reset;
  wire [63:0] regs_54_io_in;
  wire [63:0] regs_54_io_init;
  wire [63:0] regs_54_io_out;
  wire  regs_54_io_enable;
  wire  regs_55_clock;
  wire  regs_55_reset;
  wire [63:0] regs_55_io_in;
  wire [63:0] regs_55_io_init;
  wire [63:0] regs_55_io_out;
  wire  regs_55_io_enable;
  wire  regs_56_clock;
  wire  regs_56_reset;
  wire [63:0] regs_56_io_in;
  wire [63:0] regs_56_io_init;
  wire [63:0] regs_56_io_out;
  wire  regs_56_io_enable;
  wire  regs_57_clock;
  wire  regs_57_reset;
  wire [63:0] regs_57_io_in;
  wire [63:0] regs_57_io_init;
  wire [63:0] regs_57_io_out;
  wire  regs_57_io_enable;
  wire  regs_58_clock;
  wire  regs_58_reset;
  wire [63:0] regs_58_io_in;
  wire [63:0] regs_58_io_init;
  wire [63:0] regs_58_io_out;
  wire  regs_58_io_enable;
  wire  regs_59_clock;
  wire  regs_59_reset;
  wire [63:0] regs_59_io_in;
  wire [63:0] regs_59_io_init;
  wire [63:0] regs_59_io_out;
  wire  regs_59_io_enable;
  wire  regs_60_clock;
  wire  regs_60_reset;
  wire [63:0] regs_60_io_in;
  wire [63:0] regs_60_io_init;
  wire [63:0] regs_60_io_out;
  wire  regs_60_io_enable;
  wire  regs_61_clock;
  wire  regs_61_reset;
  wire [63:0] regs_61_io_in;
  wire [63:0] regs_61_io_init;
  wire [63:0] regs_61_io_out;
  wire  regs_61_io_enable;
  wire  regs_62_clock;
  wire  regs_62_reset;
  wire [63:0] regs_62_io_in;
  wire [63:0] regs_62_io_init;
  wire [63:0] regs_62_io_out;
  wire  regs_62_io_enable;
  wire  regs_63_clock;
  wire  regs_63_reset;
  wire [63:0] regs_63_io_in;
  wire [63:0] regs_63_io_init;
  wire [63:0] regs_63_io_out;
  wire  regs_63_io_enable;
  wire  regs_64_clock;
  wire  regs_64_reset;
  wire [63:0] regs_64_io_in;
  wire [63:0] regs_64_io_init;
  wire [63:0] regs_64_io_out;
  wire  regs_64_io_enable;
  wire  regs_65_clock;
  wire  regs_65_reset;
  wire [63:0] regs_65_io_in;
  wire [63:0] regs_65_io_init;
  wire [63:0] regs_65_io_out;
  wire  regs_65_io_enable;
  wire  regs_66_clock;
  wire  regs_66_reset;
  wire [63:0] regs_66_io_in;
  wire [63:0] regs_66_io_init;
  wire [63:0] regs_66_io_out;
  wire  regs_66_io_enable;
  wire  regs_67_clock;
  wire  regs_67_reset;
  wire [63:0] regs_67_io_in;
  wire [63:0] regs_67_io_init;
  wire [63:0] regs_67_io_out;
  wire  regs_67_io_enable;
  wire  regs_68_clock;
  wire  regs_68_reset;
  wire [63:0] regs_68_io_in;
  wire [63:0] regs_68_io_init;
  wire [63:0] regs_68_io_out;
  wire  regs_68_io_enable;
  wire  regs_69_clock;
  wire  regs_69_reset;
  wire [63:0] regs_69_io_in;
  wire [63:0] regs_69_io_init;
  wire [63:0] regs_69_io_out;
  wire  regs_69_io_enable;
  wire  regs_70_clock;
  wire  regs_70_reset;
  wire [63:0] regs_70_io_in;
  wire [63:0] regs_70_io_init;
  wire [63:0] regs_70_io_out;
  wire  regs_70_io_enable;
  wire  regs_71_clock;
  wire  regs_71_reset;
  wire [63:0] regs_71_io_in;
  wire [63:0] regs_71_io_init;
  wire [63:0] regs_71_io_out;
  wire  regs_71_io_enable;
  wire  regs_72_clock;
  wire  regs_72_reset;
  wire [63:0] regs_72_io_in;
  wire [63:0] regs_72_io_init;
  wire [63:0] regs_72_io_out;
  wire  regs_72_io_enable;
  wire  regs_73_clock;
  wire  regs_73_reset;
  wire [63:0] regs_73_io_in;
  wire [63:0] regs_73_io_init;
  wire [63:0] regs_73_io_out;
  wire  regs_73_io_enable;
  wire  regs_74_clock;
  wire  regs_74_reset;
  wire [63:0] regs_74_io_in;
  wire [63:0] regs_74_io_init;
  wire [63:0] regs_74_io_out;
  wire  regs_74_io_enable;
  wire  regs_75_clock;
  wire  regs_75_reset;
  wire [63:0] regs_75_io_in;
  wire [63:0] regs_75_io_init;
  wire [63:0] regs_75_io_out;
  wire  regs_75_io_enable;
  wire  regs_76_clock;
  wire  regs_76_reset;
  wire [63:0] regs_76_io_in;
  wire [63:0] regs_76_io_init;
  wire [63:0] regs_76_io_out;
  wire  regs_76_io_enable;
  wire  regs_77_clock;
  wire  regs_77_reset;
  wire [63:0] regs_77_io_in;
  wire [63:0] regs_77_io_init;
  wire [63:0] regs_77_io_out;
  wire  regs_77_io_enable;
  wire  regs_78_clock;
  wire  regs_78_reset;
  wire [63:0] regs_78_io_in;
  wire [63:0] regs_78_io_init;
  wire [63:0] regs_78_io_out;
  wire  regs_78_io_enable;
  wire  regs_79_clock;
  wire  regs_79_reset;
  wire [63:0] regs_79_io_in;
  wire [63:0] regs_79_io_init;
  wire [63:0] regs_79_io_out;
  wire  regs_79_io_enable;
  wire  regs_80_clock;
  wire  regs_80_reset;
  wire [63:0] regs_80_io_in;
  wire [63:0] regs_80_io_init;
  wire [63:0] regs_80_io_out;
  wire  regs_80_io_enable;
  wire  regs_81_clock;
  wire  regs_81_reset;
  wire [63:0] regs_81_io_in;
  wire [63:0] regs_81_io_init;
  wire [63:0] regs_81_io_out;
  wire  regs_81_io_enable;
  wire  regs_82_clock;
  wire  regs_82_reset;
  wire [63:0] regs_82_io_in;
  wire [63:0] regs_82_io_init;
  wire [63:0] regs_82_io_out;
  wire  regs_82_io_enable;
  wire  regs_83_clock;
  wire  regs_83_reset;
  wire [63:0] regs_83_io_in;
  wire [63:0] regs_83_io_init;
  wire [63:0] regs_83_io_out;
  wire  regs_83_io_enable;
  wire  regs_84_clock;
  wire  regs_84_reset;
  wire [63:0] regs_84_io_in;
  wire [63:0] regs_84_io_init;
  wire [63:0] regs_84_io_out;
  wire  regs_84_io_enable;
  wire  regs_85_clock;
  wire  regs_85_reset;
  wire [63:0] regs_85_io_in;
  wire [63:0] regs_85_io_init;
  wire [63:0] regs_85_io_out;
  wire  regs_85_io_enable;
  wire  regs_86_clock;
  wire  regs_86_reset;
  wire [63:0] regs_86_io_in;
  wire [63:0] regs_86_io_init;
  wire [63:0] regs_86_io_out;
  wire  regs_86_io_enable;
  wire  regs_87_clock;
  wire  regs_87_reset;
  wire [63:0] regs_87_io_in;
  wire [63:0] regs_87_io_init;
  wire [63:0] regs_87_io_out;
  wire  regs_87_io_enable;
  wire  regs_88_clock;
  wire  regs_88_reset;
  wire [63:0] regs_88_io_in;
  wire [63:0] regs_88_io_init;
  wire [63:0] regs_88_io_out;
  wire  regs_88_io_enable;
  wire  regs_89_clock;
  wire  regs_89_reset;
  wire [63:0] regs_89_io_in;
  wire [63:0] regs_89_io_init;
  wire [63:0] regs_89_io_out;
  wire  regs_89_io_enable;
  wire  regs_90_clock;
  wire  regs_90_reset;
  wire [63:0] regs_90_io_in;
  wire [63:0] regs_90_io_init;
  wire [63:0] regs_90_io_out;
  wire  regs_90_io_enable;
  wire  regs_91_clock;
  wire  regs_91_reset;
  wire [63:0] regs_91_io_in;
  wire [63:0] regs_91_io_init;
  wire [63:0] regs_91_io_out;
  wire  regs_91_io_enable;
  wire  regs_92_clock;
  wire  regs_92_reset;
  wire [63:0] regs_92_io_in;
  wire [63:0] regs_92_io_init;
  wire [63:0] regs_92_io_out;
  wire  regs_92_io_enable;
  wire  regs_93_clock;
  wire  regs_93_reset;
  wire [63:0] regs_93_io_in;
  wire [63:0] regs_93_io_init;
  wire [63:0] regs_93_io_out;
  wire  regs_93_io_enable;
  wire  regs_94_clock;
  wire  regs_94_reset;
  wire [63:0] regs_94_io_in;
  wire [63:0] regs_94_io_init;
  wire [63:0] regs_94_io_out;
  wire  regs_94_io_enable;
  wire  regs_95_clock;
  wire  regs_95_reset;
  wire [63:0] regs_95_io_in;
  wire [63:0] regs_95_io_init;
  wire [63:0] regs_95_io_out;
  wire  regs_95_io_enable;
  wire  regs_96_clock;
  wire  regs_96_reset;
  wire [63:0] regs_96_io_in;
  wire [63:0] regs_96_io_init;
  wire [63:0] regs_96_io_out;
  wire  regs_96_io_enable;
  wire  regs_97_clock;
  wire  regs_97_reset;
  wire [63:0] regs_97_io_in;
  wire [63:0] regs_97_io_init;
  wire [63:0] regs_97_io_out;
  wire  regs_97_io_enable;
  wire  regs_98_clock;
  wire  regs_98_reset;
  wire [63:0] regs_98_io_in;
  wire [63:0] regs_98_io_init;
  wire [63:0] regs_98_io_out;
  wire  regs_98_io_enable;
  wire  regs_99_clock;
  wire  regs_99_reset;
  wire [63:0] regs_99_io_in;
  wire [63:0] regs_99_io_init;
  wire [63:0] regs_99_io_out;
  wire  regs_99_io_enable;
  wire  regs_100_clock;
  wire  regs_100_reset;
  wire [63:0] regs_100_io_in;
  wire [63:0] regs_100_io_init;
  wire [63:0] regs_100_io_out;
  wire  regs_100_io_enable;
  wire  regs_101_clock;
  wire  regs_101_reset;
  wire [63:0] regs_101_io_in;
  wire [63:0] regs_101_io_init;
  wire [63:0] regs_101_io_out;
  wire  regs_101_io_enable;
  wire  regs_102_clock;
  wire  regs_102_reset;
  wire [63:0] regs_102_io_in;
  wire [63:0] regs_102_io_init;
  wire [63:0] regs_102_io_out;
  wire  regs_102_io_enable;
  wire  regs_103_clock;
  wire  regs_103_reset;
  wire [63:0] regs_103_io_in;
  wire [63:0] regs_103_io_init;
  wire [63:0] regs_103_io_out;
  wire  regs_103_io_enable;
  wire  regs_104_clock;
  wire  regs_104_reset;
  wire [63:0] regs_104_io_in;
  wire [63:0] regs_104_io_init;
  wire [63:0] regs_104_io_out;
  wire  regs_104_io_enable;
  wire  regs_105_clock;
  wire  regs_105_reset;
  wire [63:0] regs_105_io_in;
  wire [63:0] regs_105_io_init;
  wire [63:0] regs_105_io_out;
  wire  regs_105_io_enable;
  wire  regs_106_clock;
  wire  regs_106_reset;
  wire [63:0] regs_106_io_in;
  wire [63:0] regs_106_io_init;
  wire [63:0] regs_106_io_out;
  wire  regs_106_io_enable;
  wire  regs_107_clock;
  wire  regs_107_reset;
  wire [63:0] regs_107_io_in;
  wire [63:0] regs_107_io_init;
  wire [63:0] regs_107_io_out;
  wire  regs_107_io_enable;
  wire  regs_108_clock;
  wire  regs_108_reset;
  wire [63:0] regs_108_io_in;
  wire [63:0] regs_108_io_init;
  wire [63:0] regs_108_io_out;
  wire  regs_108_io_enable;
  wire  regs_109_clock;
  wire  regs_109_reset;
  wire [63:0] regs_109_io_in;
  wire [63:0] regs_109_io_init;
  wire [63:0] regs_109_io_out;
  wire  regs_109_io_enable;
  wire  regs_110_clock;
  wire  regs_110_reset;
  wire [63:0] regs_110_io_in;
  wire [63:0] regs_110_io_init;
  wire [63:0] regs_110_io_out;
  wire  regs_110_io_enable;
  wire  regs_111_clock;
  wire  regs_111_reset;
  wire [63:0] regs_111_io_in;
  wire [63:0] regs_111_io_init;
  wire [63:0] regs_111_io_out;
  wire  regs_111_io_enable;
  wire  regs_112_clock;
  wire  regs_112_reset;
  wire [63:0] regs_112_io_in;
  wire [63:0] regs_112_io_init;
  wire [63:0] regs_112_io_out;
  wire  regs_112_io_enable;
  wire  regs_113_clock;
  wire  regs_113_reset;
  wire [63:0] regs_113_io_in;
  wire [63:0] regs_113_io_init;
  wire [63:0] regs_113_io_out;
  wire  regs_113_io_enable;
  wire  regs_114_clock;
  wire  regs_114_reset;
  wire [63:0] regs_114_io_in;
  wire [63:0] regs_114_io_init;
  wire [63:0] regs_114_io_out;
  wire  regs_114_io_enable;
  wire  regs_115_clock;
  wire  regs_115_reset;
  wire [63:0] regs_115_io_in;
  wire [63:0] regs_115_io_init;
  wire [63:0] regs_115_io_out;
  wire  regs_115_io_enable;
  wire  regs_116_clock;
  wire  regs_116_reset;
  wire [63:0] regs_116_io_in;
  wire [63:0] regs_116_io_init;
  wire [63:0] regs_116_io_out;
  wire  regs_116_io_enable;
  wire  regs_117_clock;
  wire  regs_117_reset;
  wire [63:0] regs_117_io_in;
  wire [63:0] regs_117_io_init;
  wire [63:0] regs_117_io_out;
  wire  regs_117_io_enable;
  wire  regs_118_clock;
  wire  regs_118_reset;
  wire [63:0] regs_118_io_in;
  wire [63:0] regs_118_io_init;
  wire [63:0] regs_118_io_out;
  wire  regs_118_io_enable;
  wire  regs_119_clock;
  wire  regs_119_reset;
  wire [63:0] regs_119_io_in;
  wire [63:0] regs_119_io_init;
  wire [63:0] regs_119_io_out;
  wire  regs_119_io_enable;
  wire  regs_120_clock;
  wire  regs_120_reset;
  wire [63:0] regs_120_io_in;
  wire [63:0] regs_120_io_init;
  wire [63:0] regs_120_io_out;
  wire  regs_120_io_enable;
  wire  regs_121_clock;
  wire  regs_121_reset;
  wire [63:0] regs_121_io_in;
  wire [63:0] regs_121_io_init;
  wire [63:0] regs_121_io_out;
  wire  regs_121_io_enable;
  wire  regs_122_clock;
  wire  regs_122_reset;
  wire [63:0] regs_122_io_in;
  wire [63:0] regs_122_io_init;
  wire [63:0] regs_122_io_out;
  wire  regs_122_io_enable;
  wire  regs_123_clock;
  wire  regs_123_reset;
  wire [63:0] regs_123_io_in;
  wire [63:0] regs_123_io_init;
  wire [63:0] regs_123_io_out;
  wire  regs_123_io_enable;
  wire  regs_124_clock;
  wire  regs_124_reset;
  wire [63:0] regs_124_io_in;
  wire [63:0] regs_124_io_init;
  wire [63:0] regs_124_io_out;
  wire  regs_124_io_enable;
  wire  regs_125_clock;
  wire  regs_125_reset;
  wire [63:0] regs_125_io_in;
  wire [63:0] regs_125_io_init;
  wire [63:0] regs_125_io_out;
  wire  regs_125_io_enable;
  wire  regs_126_clock;
  wire  regs_126_reset;
  wire [63:0] regs_126_io_in;
  wire [63:0] regs_126_io_init;
  wire [63:0] regs_126_io_out;
  wire  regs_126_io_enable;
  wire  regs_127_clock;
  wire  regs_127_reset;
  wire [63:0] regs_127_io_in;
  wire [63:0] regs_127_io_init;
  wire [63:0] regs_127_io_out;
  wire  regs_127_io_enable;
  wire  regs_128_clock;
  wire  regs_128_reset;
  wire [63:0] regs_128_io_in;
  wire [63:0] regs_128_io_init;
  wire [63:0] regs_128_io_out;
  wire  regs_128_io_enable;
  wire  regs_129_clock;
  wire  regs_129_reset;
  wire [63:0] regs_129_io_in;
  wire [63:0] regs_129_io_init;
  wire [63:0] regs_129_io_out;
  wire  regs_129_io_enable;
  wire  regs_130_clock;
  wire  regs_130_reset;
  wire [63:0] regs_130_io_in;
  wire [63:0] regs_130_io_init;
  wire [63:0] regs_130_io_out;
  wire  regs_130_io_enable;
  wire  regs_131_clock;
  wire  regs_131_reset;
  wire [63:0] regs_131_io_in;
  wire [63:0] regs_131_io_init;
  wire [63:0] regs_131_io_out;
  wire  regs_131_io_enable;
  wire  regs_132_clock;
  wire  regs_132_reset;
  wire [63:0] regs_132_io_in;
  wire [63:0] regs_132_io_init;
  wire [63:0] regs_132_io_out;
  wire  regs_132_io_enable;
  wire  regs_133_clock;
  wire  regs_133_reset;
  wire [63:0] regs_133_io_in;
  wire [63:0] regs_133_io_init;
  wire [63:0] regs_133_io_out;
  wire  regs_133_io_enable;
  wire  regs_134_clock;
  wire  regs_134_reset;
  wire [63:0] regs_134_io_in;
  wire [63:0] regs_134_io_init;
  wire [63:0] regs_134_io_out;
  wire  regs_134_io_enable;
  wire  regs_135_clock;
  wire  regs_135_reset;
  wire [63:0] regs_135_io_in;
  wire [63:0] regs_135_io_init;
  wire [63:0] regs_135_io_out;
  wire  regs_135_io_enable;
  wire  regs_136_clock;
  wire  regs_136_reset;
  wire [63:0] regs_136_io_in;
  wire [63:0] regs_136_io_init;
  wire [63:0] regs_136_io_out;
  wire  regs_136_io_enable;
  wire  regs_137_clock;
  wire  regs_137_reset;
  wire [63:0] regs_137_io_in;
  wire [63:0] regs_137_io_init;
  wire [63:0] regs_137_io_out;
  wire  regs_137_io_enable;
  wire  regs_138_clock;
  wire  regs_138_reset;
  wire [63:0] regs_138_io_in;
  wire [63:0] regs_138_io_init;
  wire [63:0] regs_138_io_out;
  wire  regs_138_io_enable;
  wire  regs_139_clock;
  wire  regs_139_reset;
  wire [63:0] regs_139_io_in;
  wire [63:0] regs_139_io_init;
  wire [63:0] regs_139_io_out;
  wire  regs_139_io_enable;
  wire  regs_140_clock;
  wire  regs_140_reset;
  wire [63:0] regs_140_io_in;
  wire [63:0] regs_140_io_init;
  wire [63:0] regs_140_io_out;
  wire  regs_140_io_enable;
  wire  regs_141_clock;
  wire  regs_141_reset;
  wire [63:0] regs_141_io_in;
  wire [63:0] regs_141_io_init;
  wire [63:0] regs_141_io_out;
  wire  regs_141_io_enable;
  wire  regs_142_clock;
  wire  regs_142_reset;
  wire [63:0] regs_142_io_in;
  wire [63:0] regs_142_io_init;
  wire [63:0] regs_142_io_out;
  wire  regs_142_io_enable;
  wire  regs_143_clock;
  wire  regs_143_reset;
  wire [63:0] regs_143_io_in;
  wire [63:0] regs_143_io_init;
  wire [63:0] regs_143_io_out;
  wire  regs_143_io_enable;
  wire  regs_144_clock;
  wire  regs_144_reset;
  wire [63:0] regs_144_io_in;
  wire [63:0] regs_144_io_init;
  wire [63:0] regs_144_io_out;
  wire  regs_144_io_enable;
  wire  regs_145_clock;
  wire  regs_145_reset;
  wire [63:0] regs_145_io_in;
  wire [63:0] regs_145_io_init;
  wire [63:0] regs_145_io_out;
  wire  regs_145_io_enable;
  wire  regs_146_clock;
  wire  regs_146_reset;
  wire [63:0] regs_146_io_in;
  wire [63:0] regs_146_io_init;
  wire [63:0] regs_146_io_out;
  wire  regs_146_io_enable;
  wire  regs_147_clock;
  wire  regs_147_reset;
  wire [63:0] regs_147_io_in;
  wire [63:0] regs_147_io_init;
  wire [63:0] regs_147_io_out;
  wire  regs_147_io_enable;
  wire  regs_148_clock;
  wire  regs_148_reset;
  wire [63:0] regs_148_io_in;
  wire [63:0] regs_148_io_init;
  wire [63:0] regs_148_io_out;
  wire  regs_148_io_enable;
  wire  regs_149_clock;
  wire  regs_149_reset;
  wire [63:0] regs_149_io_in;
  wire [63:0] regs_149_io_init;
  wire [63:0] regs_149_io_out;
  wire  regs_149_io_enable;
  wire  regs_150_clock;
  wire  regs_150_reset;
  wire [63:0] regs_150_io_in;
  wire [63:0] regs_150_io_init;
  wire [63:0] regs_150_io_out;
  wire  regs_150_io_enable;
  wire  regs_151_clock;
  wire  regs_151_reset;
  wire [63:0] regs_151_io_in;
  wire [63:0] regs_151_io_init;
  wire [63:0] regs_151_io_out;
  wire  regs_151_io_enable;
  wire  regs_152_clock;
  wire  regs_152_reset;
  wire [63:0] regs_152_io_in;
  wire [63:0] regs_152_io_init;
  wire [63:0] regs_152_io_out;
  wire  regs_152_io_enable;
  wire  regs_153_clock;
  wire  regs_153_reset;
  wire [63:0] regs_153_io_in;
  wire [63:0] regs_153_io_init;
  wire [63:0] regs_153_io_out;
  wire  regs_153_io_enable;
  wire  regs_154_clock;
  wire  regs_154_reset;
  wire [63:0] regs_154_io_in;
  wire [63:0] regs_154_io_init;
  wire [63:0] regs_154_io_out;
  wire  regs_154_io_enable;
  wire  regs_155_clock;
  wire  regs_155_reset;
  wire [63:0] regs_155_io_in;
  wire [63:0] regs_155_io_init;
  wire [63:0] regs_155_io_out;
  wire  regs_155_io_enable;
  wire  regs_156_clock;
  wire  regs_156_reset;
  wire [63:0] regs_156_io_in;
  wire [63:0] regs_156_io_init;
  wire [63:0] regs_156_io_out;
  wire  regs_156_io_enable;
  wire  regs_157_clock;
  wire  regs_157_reset;
  wire [63:0] regs_157_io_in;
  wire [63:0] regs_157_io_init;
  wire [63:0] regs_157_io_out;
  wire  regs_157_io_enable;
  wire  regs_158_clock;
  wire  regs_158_reset;
  wire [63:0] regs_158_io_in;
  wire [63:0] regs_158_io_init;
  wire [63:0] regs_158_io_out;
  wire  regs_158_io_enable;
  wire  regs_159_clock;
  wire  regs_159_reset;
  wire [63:0] regs_159_io_in;
  wire [63:0] regs_159_io_init;
  wire [63:0] regs_159_io_out;
  wire  regs_159_io_enable;
  wire  regs_160_clock;
  wire  regs_160_reset;
  wire [63:0] regs_160_io_in;
  wire [63:0] regs_160_io_init;
  wire [63:0] regs_160_io_out;
  wire  regs_160_io_enable;
  wire  regs_161_clock;
  wire  regs_161_reset;
  wire [63:0] regs_161_io_in;
  wire [63:0] regs_161_io_init;
  wire [63:0] regs_161_io_out;
  wire  regs_161_io_enable;
  wire  regs_162_clock;
  wire  regs_162_reset;
  wire [63:0] regs_162_io_in;
  wire [63:0] regs_162_io_init;
  wire [63:0] regs_162_io_out;
  wire  regs_162_io_enable;
  wire  regs_163_clock;
  wire  regs_163_reset;
  wire [63:0] regs_163_io_in;
  wire [63:0] regs_163_io_init;
  wire [63:0] regs_163_io_out;
  wire  regs_163_io_enable;
  wire  regs_164_clock;
  wire  regs_164_reset;
  wire [63:0] regs_164_io_in;
  wire [63:0] regs_164_io_init;
  wire [63:0] regs_164_io_out;
  wire  regs_164_io_enable;
  wire  regs_165_clock;
  wire  regs_165_reset;
  wire [63:0] regs_165_io_in;
  wire [63:0] regs_165_io_init;
  wire [63:0] regs_165_io_out;
  wire  regs_165_io_enable;
  wire  regs_166_clock;
  wire  regs_166_reset;
  wire [63:0] regs_166_io_in;
  wire [63:0] regs_166_io_init;
  wire [63:0] regs_166_io_out;
  wire  regs_166_io_enable;
  wire  regs_167_clock;
  wire  regs_167_reset;
  wire [63:0] regs_167_io_in;
  wire [63:0] regs_167_io_init;
  wire [63:0] regs_167_io_out;
  wire  regs_167_io_enable;
  wire  regs_168_clock;
  wire  regs_168_reset;
  wire [63:0] regs_168_io_in;
  wire [63:0] regs_168_io_init;
  wire [63:0] regs_168_io_out;
  wire  regs_168_io_enable;
  wire  regs_169_clock;
  wire  regs_169_reset;
  wire [63:0] regs_169_io_in;
  wire [63:0] regs_169_io_init;
  wire [63:0] regs_169_io_out;
  wire  regs_169_io_enable;
  wire  regs_170_clock;
  wire  regs_170_reset;
  wire [63:0] regs_170_io_in;
  wire [63:0] regs_170_io_init;
  wire [63:0] regs_170_io_out;
  wire  regs_170_io_enable;
  wire  regs_171_clock;
  wire  regs_171_reset;
  wire [63:0] regs_171_io_in;
  wire [63:0] regs_171_io_init;
  wire [63:0] regs_171_io_out;
  wire  regs_171_io_enable;
  wire  regs_172_clock;
  wire  regs_172_reset;
  wire [63:0] regs_172_io_in;
  wire [63:0] regs_172_io_init;
  wire [63:0] regs_172_io_out;
  wire  regs_172_io_enable;
  wire  regs_173_clock;
  wire  regs_173_reset;
  wire [63:0] regs_173_io_in;
  wire [63:0] regs_173_io_init;
  wire [63:0] regs_173_io_out;
  wire  regs_173_io_enable;
  wire  regs_174_clock;
  wire  regs_174_reset;
  wire [63:0] regs_174_io_in;
  wire [63:0] regs_174_io_init;
  wire [63:0] regs_174_io_out;
  wire  regs_174_io_enable;
  wire  regs_175_clock;
  wire  regs_175_reset;
  wire [63:0] regs_175_io_in;
  wire [63:0] regs_175_io_init;
  wire [63:0] regs_175_io_out;
  wire  regs_175_io_enable;
  wire  regs_176_clock;
  wire  regs_176_reset;
  wire [63:0] regs_176_io_in;
  wire [63:0] regs_176_io_init;
  wire [63:0] regs_176_io_out;
  wire  regs_176_io_enable;
  wire  regs_177_clock;
  wire  regs_177_reset;
  wire [63:0] regs_177_io_in;
  wire [63:0] regs_177_io_init;
  wire [63:0] regs_177_io_out;
  wire  regs_177_io_enable;
  wire  regs_178_clock;
  wire  regs_178_reset;
  wire [63:0] regs_178_io_in;
  wire [63:0] regs_178_io_init;
  wire [63:0] regs_178_io_out;
  wire  regs_178_io_enable;
  wire  regs_179_clock;
  wire  regs_179_reset;
  wire [63:0] regs_179_io_in;
  wire [63:0] regs_179_io_init;
  wire [63:0] regs_179_io_out;
  wire  regs_179_io_enable;
  wire  regs_180_clock;
  wire  regs_180_reset;
  wire [63:0] regs_180_io_in;
  wire [63:0] regs_180_io_init;
  wire [63:0] regs_180_io_out;
  wire  regs_180_io_enable;
  wire  regs_181_clock;
  wire  regs_181_reset;
  wire [63:0] regs_181_io_in;
  wire [63:0] regs_181_io_init;
  wire [63:0] regs_181_io_out;
  wire  regs_181_io_enable;
  wire  regs_182_clock;
  wire  regs_182_reset;
  wire [63:0] regs_182_io_in;
  wire [63:0] regs_182_io_init;
  wire [63:0] regs_182_io_out;
  wire  regs_182_io_enable;
  wire  regs_183_clock;
  wire  regs_183_reset;
  wire [63:0] regs_183_io_in;
  wire [63:0] regs_183_io_init;
  wire [63:0] regs_183_io_out;
  wire  regs_183_io_enable;
  wire  regs_184_clock;
  wire  regs_184_reset;
  wire [63:0] regs_184_io_in;
  wire [63:0] regs_184_io_init;
  wire [63:0] regs_184_io_out;
  wire  regs_184_io_enable;
  wire  regs_185_clock;
  wire  regs_185_reset;
  wire [63:0] regs_185_io_in;
  wire [63:0] regs_185_io_init;
  wire [63:0] regs_185_io_out;
  wire  regs_185_io_enable;
  wire  regs_186_clock;
  wire  regs_186_reset;
  wire [63:0] regs_186_io_in;
  wire [63:0] regs_186_io_init;
  wire [63:0] regs_186_io_out;
  wire  regs_186_io_enable;
  wire  regs_187_clock;
  wire  regs_187_reset;
  wire [63:0] regs_187_io_in;
  wire [63:0] regs_187_io_init;
  wire [63:0] regs_187_io_out;
  wire  regs_187_io_enable;
  wire  regs_188_clock;
  wire  regs_188_reset;
  wire [63:0] regs_188_io_in;
  wire [63:0] regs_188_io_init;
  wire [63:0] regs_188_io_out;
  wire  regs_188_io_enable;
  wire  regs_189_clock;
  wire  regs_189_reset;
  wire [63:0] regs_189_io_in;
  wire [63:0] regs_189_io_init;
  wire [63:0] regs_189_io_out;
  wire  regs_189_io_enable;
  wire  regs_190_clock;
  wire  regs_190_reset;
  wire [63:0] regs_190_io_in;
  wire [63:0] regs_190_io_init;
  wire [63:0] regs_190_io_out;
  wire  regs_190_io_enable;
  wire  regs_191_clock;
  wire  regs_191_reset;
  wire [63:0] regs_191_io_in;
  wire [63:0] regs_191_io_init;
  wire [63:0] regs_191_io_out;
  wire  regs_191_io_enable;
  wire  regs_192_clock;
  wire  regs_192_reset;
  wire [63:0] regs_192_io_in;
  wire [63:0] regs_192_io_init;
  wire [63:0] regs_192_io_out;
  wire  regs_192_io_enable;
  wire  regs_193_clock;
  wire  regs_193_reset;
  wire [63:0] regs_193_io_in;
  wire [63:0] regs_193_io_init;
  wire [63:0] regs_193_io_out;
  wire  regs_193_io_enable;
  wire  regs_194_clock;
  wire  regs_194_reset;
  wire [63:0] regs_194_io_in;
  wire [63:0] regs_194_io_init;
  wire [63:0] regs_194_io_out;
  wire  regs_194_io_enable;
  wire  regs_195_clock;
  wire  regs_195_reset;
  wire [63:0] regs_195_io_in;
  wire [63:0] regs_195_io_init;
  wire [63:0] regs_195_io_out;
  wire  regs_195_io_enable;
  wire  regs_196_clock;
  wire  regs_196_reset;
  wire [63:0] regs_196_io_in;
  wire [63:0] regs_196_io_init;
  wire [63:0] regs_196_io_out;
  wire  regs_196_io_enable;
  wire  regs_197_clock;
  wire  regs_197_reset;
  wire [63:0] regs_197_io_in;
  wire [63:0] regs_197_io_init;
  wire [63:0] regs_197_io_out;
  wire  regs_197_io_enable;
  wire  regs_198_clock;
  wire  regs_198_reset;
  wire [63:0] regs_198_io_in;
  wire [63:0] regs_198_io_init;
  wire [63:0] regs_198_io_out;
  wire  regs_198_io_enable;
  wire  regs_199_clock;
  wire  regs_199_reset;
  wire [63:0] regs_199_io_in;
  wire [63:0] regs_199_io_init;
  wire [63:0] regs_199_io_out;
  wire  regs_199_io_enable;
  wire  regs_200_clock;
  wire  regs_200_reset;
  wire [63:0] regs_200_io_in;
  wire [63:0] regs_200_io_init;
  wire [63:0] regs_200_io_out;
  wire  regs_200_io_enable;
  wire  regs_201_clock;
  wire  regs_201_reset;
  wire [63:0] regs_201_io_in;
  wire [63:0] regs_201_io_init;
  wire [63:0] regs_201_io_out;
  wire  regs_201_io_enable;
  wire  regs_202_clock;
  wire  regs_202_reset;
  wire [63:0] regs_202_io_in;
  wire [63:0] regs_202_io_init;
  wire [63:0] regs_202_io_out;
  wire  regs_202_io_enable;
  wire  regs_203_clock;
  wire  regs_203_reset;
  wire [63:0] regs_203_io_in;
  wire [63:0] regs_203_io_init;
  wire [63:0] regs_203_io_out;
  wire  regs_203_io_enable;
  wire  regs_204_clock;
  wire  regs_204_reset;
  wire [63:0] regs_204_io_in;
  wire [63:0] regs_204_io_init;
  wire [63:0] regs_204_io_out;
  wire  regs_204_io_enable;
  wire  regs_205_clock;
  wire  regs_205_reset;
  wire [63:0] regs_205_io_in;
  wire [63:0] regs_205_io_init;
  wire [63:0] regs_205_io_out;
  wire  regs_205_io_enable;
  wire  regs_206_clock;
  wire  regs_206_reset;
  wire [63:0] regs_206_io_in;
  wire [63:0] regs_206_io_init;
  wire [63:0] regs_206_io_out;
  wire  regs_206_io_enable;
  wire  regs_207_clock;
  wire  regs_207_reset;
  wire [63:0] regs_207_io_in;
  wire [63:0] regs_207_io_init;
  wire [63:0] regs_207_io_out;
  wire  regs_207_io_enable;
  wire  regs_208_clock;
  wire  regs_208_reset;
  wire [63:0] regs_208_io_in;
  wire [63:0] regs_208_io_init;
  wire [63:0] regs_208_io_out;
  wire  regs_208_io_enable;
  wire  regs_209_clock;
  wire  regs_209_reset;
  wire [63:0] regs_209_io_in;
  wire [63:0] regs_209_io_init;
  wire [63:0] regs_209_io_out;
  wire  regs_209_io_enable;
  wire  regs_210_clock;
  wire  regs_210_reset;
  wire [63:0] regs_210_io_in;
  wire [63:0] regs_210_io_init;
  wire [63:0] regs_210_io_out;
  wire  regs_210_io_enable;
  wire  regs_211_clock;
  wire  regs_211_reset;
  wire [63:0] regs_211_io_in;
  wire [63:0] regs_211_io_init;
  wire [63:0] regs_211_io_out;
  wire  regs_211_io_enable;
  wire  regs_212_clock;
  wire  regs_212_reset;
  wire [63:0] regs_212_io_in;
  wire [63:0] regs_212_io_init;
  wire [63:0] regs_212_io_out;
  wire  regs_212_io_enable;
  wire  regs_213_clock;
  wire  regs_213_reset;
  wire [63:0] regs_213_io_in;
  wire [63:0] regs_213_io_init;
  wire [63:0] regs_213_io_out;
  wire  regs_213_io_enable;
  wire  regs_214_clock;
  wire  regs_214_reset;
  wire [63:0] regs_214_io_in;
  wire [63:0] regs_214_io_init;
  wire [63:0] regs_214_io_out;
  wire  regs_214_io_enable;
  wire  regs_215_clock;
  wire  regs_215_reset;
  wire [63:0] regs_215_io_in;
  wire [63:0] regs_215_io_init;
  wire [63:0] regs_215_io_out;
  wire  regs_215_io_enable;
  wire  regs_216_clock;
  wire  regs_216_reset;
  wire [63:0] regs_216_io_in;
  wire [63:0] regs_216_io_init;
  wire [63:0] regs_216_io_out;
  wire  regs_216_io_enable;
  wire  regs_217_clock;
  wire  regs_217_reset;
  wire [63:0] regs_217_io_in;
  wire [63:0] regs_217_io_init;
  wire [63:0] regs_217_io_out;
  wire  regs_217_io_enable;
  wire  regs_218_clock;
  wire  regs_218_reset;
  wire [63:0] regs_218_io_in;
  wire [63:0] regs_218_io_init;
  wire [63:0] regs_218_io_out;
  wire  regs_218_io_enable;
  wire  regs_219_clock;
  wire  regs_219_reset;
  wire [63:0] regs_219_io_in;
  wire [63:0] regs_219_io_init;
  wire [63:0] regs_219_io_out;
  wire  regs_219_io_enable;
  wire  regs_220_clock;
  wire  regs_220_reset;
  wire [63:0] regs_220_io_in;
  wire [63:0] regs_220_io_init;
  wire [63:0] regs_220_io_out;
  wire  regs_220_io_enable;
  wire  regs_221_clock;
  wire  regs_221_reset;
  wire [63:0] regs_221_io_in;
  wire [63:0] regs_221_io_init;
  wire [63:0] regs_221_io_out;
  wire  regs_221_io_enable;
  wire  regs_222_clock;
  wire  regs_222_reset;
  wire [63:0] regs_222_io_in;
  wire [63:0] regs_222_io_init;
  wire [63:0] regs_222_io_out;
  wire  regs_222_io_enable;
  wire  regs_223_clock;
  wire  regs_223_reset;
  wire [63:0] regs_223_io_in;
  wire [63:0] regs_223_io_init;
  wire [63:0] regs_223_io_out;
  wire  regs_223_io_enable;
  wire  regs_224_clock;
  wire  regs_224_reset;
  wire [63:0] regs_224_io_in;
  wire [63:0] regs_224_io_init;
  wire [63:0] regs_224_io_out;
  wire  regs_224_io_enable;
  wire  regs_225_clock;
  wire  regs_225_reset;
  wire [63:0] regs_225_io_in;
  wire [63:0] regs_225_io_init;
  wire [63:0] regs_225_io_out;
  wire  regs_225_io_enable;
  wire  regs_226_clock;
  wire  regs_226_reset;
  wire [63:0] regs_226_io_in;
  wire [63:0] regs_226_io_init;
  wire [63:0] regs_226_io_out;
  wire  regs_226_io_enable;
  wire  regs_227_clock;
  wire  regs_227_reset;
  wire [63:0] regs_227_io_in;
  wire [63:0] regs_227_io_init;
  wire [63:0] regs_227_io_out;
  wire  regs_227_io_enable;
  wire  regs_228_clock;
  wire  regs_228_reset;
  wire [63:0] regs_228_io_in;
  wire [63:0] regs_228_io_init;
  wire [63:0] regs_228_io_out;
  wire  regs_228_io_enable;
  wire  regs_229_clock;
  wire  regs_229_reset;
  wire [63:0] regs_229_io_in;
  wire [63:0] regs_229_io_init;
  wire [63:0] regs_229_io_out;
  wire  regs_229_io_enable;
  wire  regs_230_clock;
  wire  regs_230_reset;
  wire [63:0] regs_230_io_in;
  wire [63:0] regs_230_io_init;
  wire [63:0] regs_230_io_out;
  wire  regs_230_io_enable;
  wire  regs_231_clock;
  wire  regs_231_reset;
  wire [63:0] regs_231_io_in;
  wire [63:0] regs_231_io_init;
  wire [63:0] regs_231_io_out;
  wire  regs_231_io_enable;
  wire  regs_232_clock;
  wire  regs_232_reset;
  wire [63:0] regs_232_io_in;
  wire [63:0] regs_232_io_init;
  wire [63:0] regs_232_io_out;
  wire  regs_232_io_enable;
  wire  regs_233_clock;
  wire  regs_233_reset;
  wire [63:0] regs_233_io_in;
  wire [63:0] regs_233_io_init;
  wire [63:0] regs_233_io_out;
  wire  regs_233_io_enable;
  wire  regs_234_clock;
  wire  regs_234_reset;
  wire [63:0] regs_234_io_in;
  wire [63:0] regs_234_io_init;
  wire [63:0] regs_234_io_out;
  wire  regs_234_io_enable;
  wire  regs_235_clock;
  wire  regs_235_reset;
  wire [63:0] regs_235_io_in;
  wire [63:0] regs_235_io_init;
  wire [63:0] regs_235_io_out;
  wire  regs_235_io_enable;
  wire [63:0] rport_io_ins_0;
  wire [63:0] rport_io_ins_1;
  wire [63:0] rport_io_ins_2;
  wire [63:0] rport_io_ins_3;
  wire [63:0] rport_io_ins_4;
  wire [63:0] rport_io_ins_5;
  wire [63:0] rport_io_ins_6;
  wire [63:0] rport_io_ins_7;
  wire [63:0] rport_io_ins_8;
  wire [63:0] rport_io_ins_9;
  wire [63:0] rport_io_ins_10;
  wire [63:0] rport_io_ins_11;
  wire [63:0] rport_io_ins_12;
  wire [63:0] rport_io_ins_13;
  wire [63:0] rport_io_ins_14;
  wire [63:0] rport_io_ins_15;
  wire [63:0] rport_io_ins_16;
  wire [63:0] rport_io_ins_17;
  wire [63:0] rport_io_ins_18;
  wire [63:0] rport_io_ins_19;
  wire [63:0] rport_io_ins_20;
  wire [63:0] rport_io_ins_21;
  wire [63:0] rport_io_ins_22;
  wire [63:0] rport_io_ins_23;
  wire [63:0] rport_io_ins_24;
  wire [63:0] rport_io_ins_25;
  wire [63:0] rport_io_ins_26;
  wire [63:0] rport_io_ins_27;
  wire [63:0] rport_io_ins_28;
  wire [63:0] rport_io_ins_29;
  wire [63:0] rport_io_ins_30;
  wire [63:0] rport_io_ins_31;
  wire [63:0] rport_io_ins_32;
  wire [63:0] rport_io_ins_33;
  wire [63:0] rport_io_ins_34;
  wire [63:0] rport_io_ins_35;
  wire [63:0] rport_io_ins_36;
  wire [63:0] rport_io_ins_37;
  wire [63:0] rport_io_ins_38;
  wire [63:0] rport_io_ins_39;
  wire [63:0] rport_io_ins_40;
  wire [63:0] rport_io_ins_41;
  wire [63:0] rport_io_ins_42;
  wire [63:0] rport_io_ins_43;
  wire [63:0] rport_io_ins_44;
  wire [63:0] rport_io_ins_45;
  wire [63:0] rport_io_ins_46;
  wire [63:0] rport_io_ins_47;
  wire [63:0] rport_io_ins_48;
  wire [63:0] rport_io_ins_49;
  wire [63:0] rport_io_ins_50;
  wire [63:0] rport_io_ins_51;
  wire [63:0] rport_io_ins_52;
  wire [63:0] rport_io_ins_53;
  wire [63:0] rport_io_ins_54;
  wire [63:0] rport_io_ins_55;
  wire [63:0] rport_io_ins_56;
  wire [63:0] rport_io_ins_57;
  wire [63:0] rport_io_ins_58;
  wire [63:0] rport_io_ins_59;
  wire [63:0] rport_io_ins_60;
  wire [63:0] rport_io_ins_61;
  wire [63:0] rport_io_ins_62;
  wire [63:0] rport_io_ins_63;
  wire [63:0] rport_io_ins_64;
  wire [63:0] rport_io_ins_65;
  wire [63:0] rport_io_ins_66;
  wire [63:0] rport_io_ins_67;
  wire [63:0] rport_io_ins_68;
  wire [63:0] rport_io_ins_69;
  wire [63:0] rport_io_ins_70;
  wire [63:0] rport_io_ins_71;
  wire [63:0] rport_io_ins_72;
  wire [63:0] rport_io_ins_73;
  wire [63:0] rport_io_ins_74;
  wire [63:0] rport_io_ins_75;
  wire [63:0] rport_io_ins_76;
  wire [63:0] rport_io_ins_77;
  wire [63:0] rport_io_ins_78;
  wire [63:0] rport_io_ins_79;
  wire [63:0] rport_io_ins_80;
  wire [63:0] rport_io_ins_81;
  wire [63:0] rport_io_ins_82;
  wire [63:0] rport_io_ins_83;
  wire [63:0] rport_io_ins_84;
  wire [63:0] rport_io_ins_85;
  wire [63:0] rport_io_ins_86;
  wire [63:0] rport_io_ins_87;
  wire [63:0] rport_io_ins_88;
  wire [63:0] rport_io_ins_89;
  wire [63:0] rport_io_ins_90;
  wire [63:0] rport_io_ins_91;
  wire [63:0] rport_io_ins_92;
  wire [63:0] rport_io_ins_93;
  wire [63:0] rport_io_ins_94;
  wire [63:0] rport_io_ins_95;
  wire [63:0] rport_io_ins_96;
  wire [63:0] rport_io_ins_97;
  wire [63:0] rport_io_ins_98;
  wire [63:0] rport_io_ins_99;
  wire [63:0] rport_io_ins_100;
  wire [63:0] rport_io_ins_101;
  wire [63:0] rport_io_ins_102;
  wire [63:0] rport_io_ins_103;
  wire [63:0] rport_io_ins_104;
  wire [63:0] rport_io_ins_105;
  wire [63:0] rport_io_ins_106;
  wire [63:0] rport_io_ins_107;
  wire [63:0] rport_io_ins_108;
  wire [63:0] rport_io_ins_109;
  wire [63:0] rport_io_ins_110;
  wire [63:0] rport_io_ins_111;
  wire [63:0] rport_io_ins_112;
  wire [63:0] rport_io_ins_113;
  wire [63:0] rport_io_ins_114;
  wire [63:0] rport_io_ins_115;
  wire [63:0] rport_io_ins_116;
  wire [63:0] rport_io_ins_117;
  wire [63:0] rport_io_ins_118;
  wire [63:0] rport_io_ins_119;
  wire [63:0] rport_io_ins_120;
  wire [63:0] rport_io_ins_121;
  wire [63:0] rport_io_ins_122;
  wire [63:0] rport_io_ins_123;
  wire [63:0] rport_io_ins_124;
  wire [63:0] rport_io_ins_125;
  wire [63:0] rport_io_ins_126;
  wire [63:0] rport_io_ins_127;
  wire [63:0] rport_io_ins_128;
  wire [63:0] rport_io_ins_129;
  wire [63:0] rport_io_ins_130;
  wire [63:0] rport_io_ins_131;
  wire [63:0] rport_io_ins_132;
  wire [63:0] rport_io_ins_133;
  wire [63:0] rport_io_ins_134;
  wire [63:0] rport_io_ins_135;
  wire [63:0] rport_io_ins_136;
  wire [63:0] rport_io_ins_137;
  wire [63:0] rport_io_ins_138;
  wire [63:0] rport_io_ins_139;
  wire [63:0] rport_io_ins_140;
  wire [63:0] rport_io_ins_141;
  wire [63:0] rport_io_ins_142;
  wire [63:0] rport_io_ins_143;
  wire [63:0] rport_io_ins_144;
  wire [63:0] rport_io_ins_145;
  wire [63:0] rport_io_ins_146;
  wire [63:0] rport_io_ins_147;
  wire [63:0] rport_io_ins_148;
  wire [63:0] rport_io_ins_149;
  wire [63:0] rport_io_ins_150;
  wire [63:0] rport_io_ins_151;
  wire [63:0] rport_io_ins_152;
  wire [63:0] rport_io_ins_153;
  wire [63:0] rport_io_ins_154;
  wire [63:0] rport_io_ins_155;
  wire [63:0] rport_io_ins_156;
  wire [63:0] rport_io_ins_157;
  wire [63:0] rport_io_ins_158;
  wire [63:0] rport_io_ins_159;
  wire [63:0] rport_io_ins_160;
  wire [63:0] rport_io_ins_161;
  wire [63:0] rport_io_ins_162;
  wire [63:0] rport_io_ins_163;
  wire [63:0] rport_io_ins_164;
  wire [63:0] rport_io_ins_165;
  wire [63:0] rport_io_ins_166;
  wire [63:0] rport_io_ins_167;
  wire [63:0] rport_io_ins_168;
  wire [63:0] rport_io_ins_169;
  wire [63:0] rport_io_ins_170;
  wire [63:0] rport_io_ins_171;
  wire [63:0] rport_io_ins_172;
  wire [63:0] rport_io_ins_173;
  wire [63:0] rport_io_ins_174;
  wire [63:0] rport_io_ins_175;
  wire [63:0] rport_io_ins_176;
  wire [63:0] rport_io_ins_177;
  wire [63:0] rport_io_ins_178;
  wire [63:0] rport_io_ins_179;
  wire [63:0] rport_io_ins_180;
  wire [63:0] rport_io_ins_181;
  wire [63:0] rport_io_ins_182;
  wire [63:0] rport_io_ins_183;
  wire [63:0] rport_io_ins_184;
  wire [63:0] rport_io_ins_185;
  wire [63:0] rport_io_ins_186;
  wire [63:0] rport_io_ins_187;
  wire [63:0] rport_io_ins_188;
  wire [63:0] rport_io_ins_189;
  wire [63:0] rport_io_ins_190;
  wire [63:0] rport_io_ins_191;
  wire [63:0] rport_io_ins_192;
  wire [63:0] rport_io_ins_193;
  wire [63:0] rport_io_ins_194;
  wire [63:0] rport_io_ins_195;
  wire [63:0] rport_io_ins_196;
  wire [63:0] rport_io_ins_197;
  wire [63:0] rport_io_ins_198;
  wire [63:0] rport_io_ins_199;
  wire [63:0] rport_io_ins_200;
  wire [63:0] rport_io_ins_201;
  wire [63:0] rport_io_ins_202;
  wire [63:0] rport_io_ins_203;
  wire [63:0] rport_io_ins_204;
  wire [63:0] rport_io_ins_205;
  wire [63:0] rport_io_ins_206;
  wire [63:0] rport_io_ins_207;
  wire [63:0] rport_io_ins_208;
  wire [63:0] rport_io_ins_209;
  wire [63:0] rport_io_ins_210;
  wire [63:0] rport_io_ins_211;
  wire [63:0] rport_io_ins_212;
  wire [63:0] rport_io_ins_213;
  wire [63:0] rport_io_ins_214;
  wire [63:0] rport_io_ins_215;
  wire [63:0] rport_io_ins_216;
  wire [63:0] rport_io_ins_217;
  wire [63:0] rport_io_ins_218;
  wire [63:0] rport_io_ins_219;
  wire [63:0] rport_io_ins_220;
  wire [63:0] rport_io_ins_221;
  wire [63:0] rport_io_ins_222;
  wire [63:0] rport_io_ins_223;
  wire [63:0] rport_io_ins_224;
  wire [63:0] rport_io_ins_225;
  wire [63:0] rport_io_ins_226;
  wire [63:0] rport_io_ins_227;
  wire [63:0] rport_io_ins_228;
  wire [63:0] rport_io_ins_229;
  wire [63:0] rport_io_ins_230;
  wire [63:0] rport_io_ins_231;
  wire [63:0] rport_io_ins_232;
  wire [63:0] rport_io_ins_233;
  wire [63:0] rport_io_ins_234;
  wire [63:0] rport_io_ins_235;
  wire [7:0] rport_io_sel;
  wire [63:0] rport_io_out;
  wire [63:0] regOuts_0;
  wire [63:0] regOuts_1;
  wire [63:0] regOuts_2;
  wire [63:0] regOuts_3;
  wire [63:0] regOuts_4;
  wire [63:0] regOuts_5;
  wire [63:0] regOuts_6;
  wire [63:0] regOuts_7;
  wire [63:0] regOuts_8;
  wire [63:0] regOuts_9;
  wire [63:0] regOuts_10;
  wire [63:0] regOuts_11;
  wire [63:0] regOuts_12;
  wire [63:0] regOuts_13;
  wire [63:0] regOuts_14;
  wire [63:0] regOuts_15;
  wire [63:0] regOuts_16;
  wire [63:0] regOuts_17;
  wire [63:0] regOuts_18;
  wire [63:0] regOuts_19;
  wire [63:0] regOuts_20;
  wire [63:0] regOuts_21;
  wire [63:0] regOuts_22;
  wire [63:0] regOuts_23;
  wire [63:0] regOuts_24;
  wire [63:0] regOuts_25;
  wire [63:0] regOuts_26;
  wire [63:0] regOuts_27;
  wire [63:0] regOuts_28;
  wire [63:0] regOuts_29;
  wire [63:0] regOuts_30;
  wire [63:0] regOuts_31;
  wire [63:0] regOuts_32;
  wire [63:0] regOuts_33;
  wire [63:0] regOuts_34;
  wire [63:0] regOuts_35;
  wire [63:0] regOuts_36;
  wire [63:0] regOuts_37;
  wire [63:0] regOuts_38;
  wire [63:0] regOuts_39;
  wire [63:0] regOuts_40;
  wire [63:0] regOuts_41;
  wire [63:0] regOuts_42;
  wire [63:0] regOuts_43;
  wire [63:0] regOuts_44;
  wire [63:0] regOuts_45;
  wire [63:0] regOuts_46;
  wire [63:0] regOuts_47;
  wire [63:0] regOuts_48;
  wire [63:0] regOuts_49;
  wire [63:0] regOuts_50;
  wire [63:0] regOuts_51;
  wire [63:0] regOuts_52;
  wire [63:0] regOuts_53;
  wire [63:0] regOuts_54;
  wire [63:0] regOuts_55;
  wire [63:0] regOuts_56;
  wire [63:0] regOuts_57;
  wire [63:0] regOuts_58;
  wire [63:0] regOuts_59;
  wire [63:0] regOuts_60;
  wire [63:0] regOuts_61;
  wire [63:0] regOuts_62;
  wire [63:0] regOuts_63;
  wire [63:0] regOuts_64;
  wire [63:0] regOuts_65;
  wire [63:0] regOuts_66;
  wire [63:0] regOuts_67;
  wire [63:0] regOuts_68;
  wire [63:0] regOuts_69;
  wire [63:0] regOuts_70;
  wire [63:0] regOuts_71;
  wire [63:0] regOuts_72;
  wire [63:0] regOuts_73;
  wire [63:0] regOuts_74;
  wire [63:0] regOuts_75;
  wire [63:0] regOuts_76;
  wire [63:0] regOuts_77;
  wire [63:0] regOuts_78;
  wire [63:0] regOuts_79;
  wire [63:0] regOuts_80;
  wire [63:0] regOuts_81;
  wire [63:0] regOuts_82;
  wire [63:0] regOuts_83;
  wire [63:0] regOuts_84;
  wire [63:0] regOuts_85;
  wire [63:0] regOuts_86;
  wire [63:0] regOuts_87;
  wire [63:0] regOuts_88;
  wire [63:0] regOuts_89;
  wire [63:0] regOuts_90;
  wire [63:0] regOuts_91;
  wire [63:0] regOuts_92;
  wire [63:0] regOuts_93;
  wire [63:0] regOuts_94;
  wire [63:0] regOuts_95;
  wire [63:0] regOuts_96;
  wire [63:0] regOuts_97;
  wire [63:0] regOuts_98;
  wire [63:0] regOuts_99;
  wire [63:0] regOuts_100;
  wire [63:0] regOuts_101;
  wire [63:0] regOuts_102;
  wire [63:0] regOuts_103;
  wire [63:0] regOuts_104;
  wire [63:0] regOuts_105;
  wire [63:0] regOuts_106;
  wire [63:0] regOuts_107;
  wire [63:0] regOuts_108;
  wire [63:0] regOuts_109;
  wire [63:0] regOuts_110;
  wire [63:0] regOuts_111;
  wire [63:0] regOuts_112;
  wire [63:0] regOuts_113;
  wire [63:0] regOuts_114;
  wire [63:0] regOuts_115;
  wire [63:0] regOuts_116;
  wire [63:0] regOuts_117;
  wire [63:0] regOuts_118;
  wire [63:0] regOuts_119;
  wire [63:0] regOuts_120;
  wire [63:0] regOuts_121;
  wire [63:0] regOuts_122;
  wire [63:0] regOuts_123;
  wire [63:0] regOuts_124;
  wire [63:0] regOuts_125;
  wire [63:0] regOuts_126;
  wire [63:0] regOuts_127;
  wire [63:0] regOuts_128;
  wire [63:0] regOuts_129;
  wire [63:0] regOuts_130;
  wire [63:0] regOuts_131;
  wire [63:0] regOuts_132;
  wire [63:0] regOuts_133;
  wire [63:0] regOuts_134;
  wire [63:0] regOuts_135;
  wire [63:0] regOuts_136;
  wire [63:0] regOuts_137;
  wire [63:0] regOuts_138;
  wire [63:0] regOuts_139;
  wire [63:0] regOuts_140;
  wire [63:0] regOuts_141;
  wire [63:0] regOuts_142;
  wire [63:0] regOuts_143;
  wire [63:0] regOuts_144;
  wire [63:0] regOuts_145;
  wire [63:0] regOuts_146;
  wire [63:0] regOuts_147;
  wire [63:0] regOuts_148;
  wire [63:0] regOuts_149;
  wire [63:0] regOuts_150;
  wire [63:0] regOuts_151;
  wire [63:0] regOuts_152;
  wire [63:0] regOuts_153;
  wire [63:0] regOuts_154;
  wire [63:0] regOuts_155;
  wire [63:0] regOuts_156;
  wire [63:0] regOuts_157;
  wire [63:0] regOuts_158;
  wire [63:0] regOuts_159;
  wire [63:0] regOuts_160;
  wire [63:0] regOuts_161;
  wire [63:0] regOuts_162;
  wire [63:0] regOuts_163;
  wire [63:0] regOuts_164;
  wire [63:0] regOuts_165;
  wire [63:0] regOuts_166;
  wire [63:0] regOuts_167;
  wire [63:0] regOuts_168;
  wire [63:0] regOuts_169;
  wire [63:0] regOuts_170;
  wire [63:0] regOuts_171;
  wire [63:0] regOuts_172;
  wire [63:0] regOuts_173;
  wire [63:0] regOuts_174;
  wire [63:0] regOuts_175;
  wire [63:0] regOuts_176;
  wire [63:0] regOuts_177;
  wire [63:0] regOuts_178;
  wire [63:0] regOuts_179;
  wire [63:0] regOuts_180;
  wire [63:0] regOuts_181;
  wire [63:0] regOuts_182;
  wire [63:0] regOuts_183;
  wire [63:0] regOuts_184;
  wire [63:0] regOuts_185;
  wire [63:0] regOuts_186;
  wire [63:0] regOuts_187;
  wire [63:0] regOuts_188;
  wire [63:0] regOuts_189;
  wire [63:0] regOuts_190;
  wire [63:0] regOuts_191;
  wire [63:0] regOuts_192;
  wire [63:0] regOuts_193;
  wire [63:0] regOuts_194;
  wire [63:0] regOuts_195;
  wire [63:0] regOuts_196;
  wire [63:0] regOuts_197;
  wire [63:0] regOuts_198;
  wire [63:0] regOuts_199;
  wire [63:0] regOuts_200;
  wire [63:0] regOuts_201;
  wire [63:0] regOuts_202;
  wire [63:0] regOuts_203;
  wire [63:0] regOuts_204;
  wire [63:0] regOuts_205;
  wire [63:0] regOuts_206;
  wire [63:0] regOuts_207;
  wire [63:0] regOuts_208;
  wire [63:0] regOuts_209;
  wire [63:0] regOuts_210;
  wire [63:0] regOuts_211;
  wire [63:0] regOuts_212;
  wire [63:0] regOuts_213;
  wire [63:0] regOuts_214;
  wire [63:0] regOuts_215;
  wire [63:0] regOuts_216;
  wire [63:0] regOuts_217;
  wire [63:0] regOuts_218;
  wire [63:0] regOuts_219;
  wire [63:0] regOuts_220;
  wire [63:0] regOuts_221;
  wire [63:0] regOuts_222;
  wire [63:0] regOuts_223;
  wire [63:0] regOuts_224;
  wire [63:0] regOuts_225;
  wire [63:0] regOuts_226;
  wire [63:0] regOuts_227;
  wire [63:0] regOuts_228;
  wire [63:0] regOuts_229;
  wire [63:0] regOuts_230;
  wire [63:0] regOuts_231;
  wire [63:0] regOuts_232;
  wire [63:0] regOuts_233;
  wire [63:0] regOuts_234;
  wire [63:0] regOuts_235;
  wire [63:0] _T_2390_0;
  wire [63:0] _T_2390_1;
  wire [63:0] _T_2390_2;
  FF_1160 regs_0 (
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_init(regs_0_io_init),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FF_1160 regs_1 (
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_init(regs_1_io_init),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FF_1160 regs_2 (
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_init(regs_2_io_init),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FF_1160 regs_3 (
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_init(regs_3_io_init),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FF_1160 regs_4 (
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_init(regs_4_io_init),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FF_1160 regs_5 (
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_init(regs_5_io_init),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FF_1160 regs_6 (
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_init(regs_6_io_init),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FF_1160 regs_7 (
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_init(regs_7_io_init),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FF_1160 regs_8 (
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_init(regs_8_io_init),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FF_1160 regs_9 (
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_init(regs_9_io_init),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FF_1160 regs_10 (
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_init(regs_10_io_init),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FF_1160 regs_11 (
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_init(regs_11_io_init),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FF_1160 regs_12 (
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_init(regs_12_io_init),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FF_1160 regs_13 (
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_init(regs_13_io_init),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FF_1160 regs_14 (
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_init(regs_14_io_init),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FF_1160 regs_15 (
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_init(regs_15_io_init),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FF_1160 regs_16 (
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_init(regs_16_io_init),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FF_1160 regs_17 (
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_init(regs_17_io_init),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FF_1160 regs_18 (
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_init(regs_18_io_init),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FF_1160 regs_19 (
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_init(regs_19_io_init),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FF_1160 regs_20 (
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_init(regs_20_io_init),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FF_1160 regs_21 (
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_init(regs_21_io_init),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FF_1160 regs_22 (
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_init(regs_22_io_init),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FF_1160 regs_23 (
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_init(regs_23_io_init),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FF_1160 regs_24 (
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_init(regs_24_io_init),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FF_1160 regs_25 (
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_init(regs_25_io_init),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FF_1160 regs_26 (
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_init(regs_26_io_init),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FF_1160 regs_27 (
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_init(regs_27_io_init),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FF_1160 regs_28 (
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_init(regs_28_io_init),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FF_1160 regs_29 (
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_init(regs_29_io_init),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FF_1160 regs_30 (
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_init(regs_30_io_init),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FF_1160 regs_31 (
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_init(regs_31_io_init),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FF_1160 regs_32 (
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_init(regs_32_io_init),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FF_1160 regs_33 (
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_init(regs_33_io_init),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FF_1160 regs_34 (
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_init(regs_34_io_init),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FF_1160 regs_35 (
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_init(regs_35_io_init),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FF_1160 regs_36 (
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_init(regs_36_io_init),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FF_1160 regs_37 (
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_init(regs_37_io_init),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FF_1160 regs_38 (
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_init(regs_38_io_init),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FF_1160 regs_39 (
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_init(regs_39_io_init),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FF_1160 regs_40 (
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_init(regs_40_io_init),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FF_1160 regs_41 (
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_init(regs_41_io_init),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FF_1160 regs_42 (
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_init(regs_42_io_init),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FF_1160 regs_43 (
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_init(regs_43_io_init),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FF_1160 regs_44 (
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_init(regs_44_io_init),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FF_1160 regs_45 (
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_init(regs_45_io_init),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FF_1160 regs_46 (
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_init(regs_46_io_init),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FF_1160 regs_47 (
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_init(regs_47_io_init),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FF_1160 regs_48 (
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_init(regs_48_io_init),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FF_1160 regs_49 (
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_init(regs_49_io_init),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FF_1160 regs_50 (
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_init(regs_50_io_init),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FF_1160 regs_51 (
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_init(regs_51_io_init),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FF_1160 regs_52 (
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_init(regs_52_io_init),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FF_1160 regs_53 (
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_init(regs_53_io_init),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FF_1160 regs_54 (
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_init(regs_54_io_init),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FF_1160 regs_55 (
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_init(regs_55_io_init),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FF_1160 regs_56 (
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_init(regs_56_io_init),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FF_1160 regs_57 (
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_init(regs_57_io_init),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FF_1160 regs_58 (
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_init(regs_58_io_init),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FF_1160 regs_59 (
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_init(regs_59_io_init),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FF_1160 regs_60 (
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_init(regs_60_io_init),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FF_1160 regs_61 (
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_init(regs_61_io_init),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FF_1160 regs_62 (
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_init(regs_62_io_init),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FF_1160 regs_63 (
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_init(regs_63_io_init),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FF_1160 regs_64 (
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_init(regs_64_io_init),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FF_1160 regs_65 (
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_init(regs_65_io_init),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FF_1160 regs_66 (
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_init(regs_66_io_init),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FF_1160 regs_67 (
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_init(regs_67_io_init),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FF_1160 regs_68 (
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_init(regs_68_io_init),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FF_1160 regs_69 (
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_init(regs_69_io_init),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FF_1160 regs_70 (
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_init(regs_70_io_init),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FF_1160 regs_71 (
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_init(regs_71_io_init),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FF_1160 regs_72 (
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_init(regs_72_io_init),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FF_1160 regs_73 (
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_init(regs_73_io_init),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FF_1160 regs_74 (
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_init(regs_74_io_init),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FF_1160 regs_75 (
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_init(regs_75_io_init),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FF_1160 regs_76 (
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_init(regs_76_io_init),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FF_1160 regs_77 (
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_init(regs_77_io_init),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FF_1160 regs_78 (
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_init(regs_78_io_init),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FF_1160 regs_79 (
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_init(regs_79_io_init),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FF_1160 regs_80 (
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_init(regs_80_io_init),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FF_1160 regs_81 (
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_init(regs_81_io_init),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FF_1160 regs_82 (
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_init(regs_82_io_init),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FF_1160 regs_83 (
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_init(regs_83_io_init),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FF_1160 regs_84 (
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_init(regs_84_io_init),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FF_1160 regs_85 (
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_init(regs_85_io_init),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FF_1160 regs_86 (
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_init(regs_86_io_init),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FF_1160 regs_87 (
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_init(regs_87_io_init),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FF_1160 regs_88 (
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_init(regs_88_io_init),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FF_1160 regs_89 (
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_init(regs_89_io_init),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FF_1160 regs_90 (
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_init(regs_90_io_init),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FF_1160 regs_91 (
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_init(regs_91_io_init),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FF_1160 regs_92 (
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_init(regs_92_io_init),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FF_1160 regs_93 (
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_init(regs_93_io_init),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FF_1160 regs_94 (
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_init(regs_94_io_init),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FF_1160 regs_95 (
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_init(regs_95_io_init),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FF_1160 regs_96 (
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_init(regs_96_io_init),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FF_1160 regs_97 (
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_init(regs_97_io_init),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FF_1160 regs_98 (
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_init(regs_98_io_init),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FF_1160 regs_99 (
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_init(regs_99_io_init),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FF_1160 regs_100 (
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_init(regs_100_io_init),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FF_1160 regs_101 (
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_init(regs_101_io_init),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FF_1160 regs_102 (
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_init(regs_102_io_init),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FF_1160 regs_103 (
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_init(regs_103_io_init),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FF_1160 regs_104 (
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_init(regs_104_io_init),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FF_1160 regs_105 (
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_init(regs_105_io_init),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FF_1160 regs_106 (
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_init(regs_106_io_init),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FF_1160 regs_107 (
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_init(regs_107_io_init),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FF_1160 regs_108 (
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_init(regs_108_io_init),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FF_1160 regs_109 (
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_init(regs_109_io_init),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FF_1160 regs_110 (
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_init(regs_110_io_init),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FF_1160 regs_111 (
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_init(regs_111_io_init),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FF_1160 regs_112 (
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_init(regs_112_io_init),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FF_1160 regs_113 (
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_init(regs_113_io_init),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FF_1160 regs_114 (
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_init(regs_114_io_init),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FF_1160 regs_115 (
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_init(regs_115_io_init),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FF_1160 regs_116 (
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_init(regs_116_io_init),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FF_1160 regs_117 (
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_init(regs_117_io_init),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FF_1160 regs_118 (
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_init(regs_118_io_init),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FF_1160 regs_119 (
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_init(regs_119_io_init),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FF_1160 regs_120 (
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_init(regs_120_io_init),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FF_1160 regs_121 (
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_init(regs_121_io_init),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FF_1160 regs_122 (
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_init(regs_122_io_init),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FF_1160 regs_123 (
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_init(regs_123_io_init),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FF_1160 regs_124 (
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_init(regs_124_io_init),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FF_1160 regs_125 (
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_init(regs_125_io_init),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FF_1160 regs_126 (
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_init(regs_126_io_init),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FF_1160 regs_127 (
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_init(regs_127_io_init),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FF_1160 regs_128 (
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_init(regs_128_io_init),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FF_1160 regs_129 (
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_init(regs_129_io_init),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FF_1160 regs_130 (
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_init(regs_130_io_init),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FF_1160 regs_131 (
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_init(regs_131_io_init),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FF_1160 regs_132 (
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_init(regs_132_io_init),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FF_1160 regs_133 (
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_init(regs_133_io_init),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FF_1160 regs_134 (
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_init(regs_134_io_init),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FF_1160 regs_135 (
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_init(regs_135_io_init),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FF_1160 regs_136 (
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_init(regs_136_io_init),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FF_1160 regs_137 (
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_init(regs_137_io_init),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FF_1160 regs_138 (
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_init(regs_138_io_init),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FF_1160 regs_139 (
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_init(regs_139_io_init),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FF_1160 regs_140 (
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_init(regs_140_io_init),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FF_1160 regs_141 (
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_init(regs_141_io_init),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FF_1160 regs_142 (
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_init(regs_142_io_init),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FF_1160 regs_143 (
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_init(regs_143_io_init),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FF_1160 regs_144 (
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_init(regs_144_io_init),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FF_1160 regs_145 (
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_init(regs_145_io_init),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FF_1160 regs_146 (
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_init(regs_146_io_init),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FF_1160 regs_147 (
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_init(regs_147_io_init),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FF_1160 regs_148 (
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_init(regs_148_io_init),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FF_1160 regs_149 (
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_init(regs_149_io_init),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FF_1160 regs_150 (
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_init(regs_150_io_init),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FF_1160 regs_151 (
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_init(regs_151_io_init),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FF_1160 regs_152 (
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_init(regs_152_io_init),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FF_1160 regs_153 (
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_init(regs_153_io_init),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FF_1160 regs_154 (
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_init(regs_154_io_init),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FF_1160 regs_155 (
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_init(regs_155_io_init),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FF_1160 regs_156 (
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_init(regs_156_io_init),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FF_1160 regs_157 (
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_init(regs_157_io_init),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FF_1160 regs_158 (
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_init(regs_158_io_init),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FF_1160 regs_159 (
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_init(regs_159_io_init),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FF_1160 regs_160 (
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_init(regs_160_io_init),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FF_1160 regs_161 (
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_init(regs_161_io_init),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FF_1160 regs_162 (
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_init(regs_162_io_init),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FF_1160 regs_163 (
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_init(regs_163_io_init),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FF_1160 regs_164 (
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_init(regs_164_io_init),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FF_1160 regs_165 (
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_init(regs_165_io_init),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FF_1160 regs_166 (
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_init(regs_166_io_init),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FF_1160 regs_167 (
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_init(regs_167_io_init),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FF_1160 regs_168 (
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_init(regs_168_io_init),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FF_1160 regs_169 (
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_init(regs_169_io_init),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FF_1160 regs_170 (
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_init(regs_170_io_init),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FF_1160 regs_171 (
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_init(regs_171_io_init),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FF_1160 regs_172 (
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_init(regs_172_io_init),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FF_1160 regs_173 (
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_init(regs_173_io_init),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FF_1160 regs_174 (
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_init(regs_174_io_init),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FF_1160 regs_175 (
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_init(regs_175_io_init),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FF_1160 regs_176 (
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_init(regs_176_io_init),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FF_1160 regs_177 (
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_init(regs_177_io_init),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FF_1160 regs_178 (
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_init(regs_178_io_init),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FF_1160 regs_179 (
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_init(regs_179_io_init),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FF_1160 regs_180 (
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_init(regs_180_io_init),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FF_1160 regs_181 (
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_init(regs_181_io_init),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FF_1160 regs_182 (
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_init(regs_182_io_init),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FF_1160 regs_183 (
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_init(regs_183_io_init),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FF_1160 regs_184 (
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_init(regs_184_io_init),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FF_1160 regs_185 (
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_init(regs_185_io_init),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FF_1160 regs_186 (
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_init(regs_186_io_init),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FF_1160 regs_187 (
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_init(regs_187_io_init),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FF_1160 regs_188 (
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_init(regs_188_io_init),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FF_1160 regs_189 (
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_init(regs_189_io_init),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FF_1160 regs_190 (
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_init(regs_190_io_init),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FF_1160 regs_191 (
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_init(regs_191_io_init),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FF_1160 regs_192 (
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_init(regs_192_io_init),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FF_1160 regs_193 (
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_init(regs_193_io_init),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FF_1160 regs_194 (
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_init(regs_194_io_init),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FF_1160 regs_195 (
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_init(regs_195_io_init),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FF_1160 regs_196 (
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_init(regs_196_io_init),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FF_1160 regs_197 (
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_init(regs_197_io_init),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FF_1160 regs_198 (
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_init(regs_198_io_init),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FF_1160 regs_199 (
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_init(regs_199_io_init),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FF_1160 regs_200 (
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_init(regs_200_io_init),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FF_1160 regs_201 (
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_init(regs_201_io_init),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FF_1160 regs_202 (
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_init(regs_202_io_init),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FF_1160 regs_203 (
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_init(regs_203_io_init),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FF_1160 regs_204 (
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_init(regs_204_io_init),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FF_1160 regs_205 (
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_init(regs_205_io_init),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FF_1160 regs_206 (
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_init(regs_206_io_init),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FF_1160 regs_207 (
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_init(regs_207_io_init),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FF_1160 regs_208 (
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_init(regs_208_io_init),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FF_1160 regs_209 (
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_init(regs_209_io_init),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FF_1160 regs_210 (
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_init(regs_210_io_init),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FF_1160 regs_211 (
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_init(regs_211_io_init),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FF_1160 regs_212 (
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_init(regs_212_io_init),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FF_1160 regs_213 (
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_init(regs_213_io_init),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FF_1160 regs_214 (
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_init(regs_214_io_init),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FF_1160 regs_215 (
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_init(regs_215_io_init),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FF_1160 regs_216 (
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_init(regs_216_io_init),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FF_1160 regs_217 (
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_init(regs_217_io_init),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FF_1160 regs_218 (
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_init(regs_218_io_init),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FF_1160 regs_219 (
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_init(regs_219_io_init),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FF_1160 regs_220 (
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_init(regs_220_io_init),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FF_1160 regs_221 (
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_init(regs_221_io_init),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FF_1160 regs_222 (
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_init(regs_222_io_init),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FF_1160 regs_223 (
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_init(regs_223_io_init),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FF_1160 regs_224 (
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_init(regs_224_io_init),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FF_1160 regs_225 (
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_init(regs_225_io_init),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FF_1160 regs_226 (
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_init(regs_226_io_init),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FF_1160 regs_227 (
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_init(regs_227_io_init),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FF_1160 regs_228 (
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_init(regs_228_io_init),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FF_1160 regs_229 (
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_init(regs_229_io_init),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FF_1160 regs_230 (
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_init(regs_230_io_init),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FF_1160 regs_231 (
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_init(regs_231_io_init),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FF_1160 regs_232 (
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_init(regs_232_io_init),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FF_1160 regs_233 (
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_init(regs_233_io_init),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FF_1160 regs_234 (
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_init(regs_234_io_init),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FF_1160 regs_235 (
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_init(regs_235_io_init),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  MuxN_6 rport (
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_731 = io_waddr == 8'h0;
  assign _T_732 = io_wen & _T_731;
  assign _T_735 = io_waddr == 8'h1;
  assign _T_736 = io_wen & _T_735;
  assign _T_740 = _T_736 ? _T_736 : io_argOuts_0_valid;
  assign _T_744 = _T_736 ? io_wdata : io_argOuts_0_bits;
  assign _T_747 = io_waddr == 8'h2;
  assign _T_748 = io_wen & _T_747;
  assign _T_751 = io_waddr == 8'h3;
  assign _T_752 = io_wen & _T_751;
  assign _T_753 = io_argOuts_1_valid | _T_752;
  assign _T_754 = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata;
  assign io_rdata = rport_io_out;
  assign io_argIns_0 = _T_2390_0;
  assign io_argIns_1 = _T_2390_1;
  assign io_argIns_2 = _T_2390_2;
  assign regs_0_io_in = io_wdata;
  assign regs_0_io_init = 64'h0;
  assign regs_0_io_enable = _T_732;
  assign regs_0_clock = clock;
  assign regs_0_reset = reset;
  assign regs_1_io_in = _T_744;
  assign regs_1_io_init = 64'h0;
  assign regs_1_io_enable = _T_740;
  assign regs_1_clock = clock;
  assign regs_1_reset = reset;
  assign regs_2_io_in = io_wdata;
  assign regs_2_io_init = 64'h0;
  assign regs_2_io_enable = _T_748;
  assign regs_2_clock = clock;
  assign regs_2_reset = reset;
  assign regs_3_io_in = _T_754;
  assign regs_3_io_init = 64'h0;
  assign regs_3_io_enable = _T_753;
  assign regs_3_clock = clock;
  assign regs_3_reset = reset;
  assign regs_4_io_in = io_argOuts_2_bits;
  assign regs_4_io_init = 64'h0;
  assign regs_4_io_enable = 1'h1;
  assign regs_4_clock = clock;
  assign regs_4_reset = reset;
  assign regs_5_io_in = io_argOuts_3_bits;
  assign regs_5_io_init = 64'h0;
  assign regs_5_io_enable = 1'h1;
  assign regs_5_clock = clock;
  assign regs_5_reset = reset;
  assign regs_6_io_in = io_argOuts_4_bits;
  assign regs_6_io_init = 64'h0;
  assign regs_6_io_enable = 1'h1;
  assign regs_6_clock = clock;
  assign regs_6_reset = reset;
  assign regs_7_io_in = io_argOuts_5_bits;
  assign regs_7_io_init = 64'h0;
  assign regs_7_io_enable = 1'h1;
  assign regs_7_clock = clock;
  assign regs_7_reset = reset;
  assign regs_8_io_in = io_argOuts_6_bits;
  assign regs_8_io_init = 64'h0;
  assign regs_8_io_enable = 1'h1;
  assign regs_8_clock = clock;
  assign regs_8_reset = reset;
  assign regs_9_io_in = io_argOuts_7_bits;
  assign regs_9_io_init = 64'h0;
  assign regs_9_io_enable = 1'h1;
  assign regs_9_clock = clock;
  assign regs_9_reset = reset;
  assign regs_10_io_in = io_argOuts_8_bits;
  assign regs_10_io_init = 64'h0;
  assign regs_10_io_enable = 1'h1;
  assign regs_10_clock = clock;
  assign regs_10_reset = reset;
  assign regs_11_io_in = io_argOuts_9_bits;
  assign regs_11_io_init = 64'h0;
  assign regs_11_io_enable = 1'h1;
  assign regs_11_clock = clock;
  assign regs_11_reset = reset;
  assign regs_12_io_in = io_argOuts_10_bits;
  assign regs_12_io_init = 64'h0;
  assign regs_12_io_enable = 1'h1;
  assign regs_12_clock = clock;
  assign regs_12_reset = reset;
  assign regs_13_io_in = io_argOuts_11_bits;
  assign regs_13_io_init = 64'h0;
  assign regs_13_io_enable = 1'h1;
  assign regs_13_clock = clock;
  assign regs_13_reset = reset;
  assign regs_14_io_in = io_argOuts_12_bits;
  assign regs_14_io_init = 64'h0;
  assign regs_14_io_enable = 1'h1;
  assign regs_14_clock = clock;
  assign regs_14_reset = reset;
  assign regs_15_io_in = io_argOuts_13_bits;
  assign regs_15_io_init = 64'h0;
  assign regs_15_io_enable = 1'h1;
  assign regs_15_clock = clock;
  assign regs_15_reset = reset;
  assign regs_16_io_in = io_argOuts_14_bits;
  assign regs_16_io_init = 64'h0;
  assign regs_16_io_enable = 1'h1;
  assign regs_16_clock = clock;
  assign regs_16_reset = reset;
  assign regs_17_io_in = io_argOuts_15_bits;
  assign regs_17_io_init = 64'h0;
  assign regs_17_io_enable = 1'h1;
  assign regs_17_clock = clock;
  assign regs_17_reset = reset;
  assign regs_18_io_in = io_argOuts_16_bits;
  assign regs_18_io_init = 64'h0;
  assign regs_18_io_enable = 1'h1;
  assign regs_18_clock = clock;
  assign regs_18_reset = reset;
  assign regs_19_io_in = io_argOuts_17_bits;
  assign regs_19_io_init = 64'h0;
  assign regs_19_io_enable = 1'h1;
  assign regs_19_clock = clock;
  assign regs_19_reset = reset;
  assign regs_20_io_in = io_argOuts_18_bits;
  assign regs_20_io_init = 64'h0;
  assign regs_20_io_enable = 1'h1;
  assign regs_20_clock = clock;
  assign regs_20_reset = reset;
  assign regs_21_io_in = io_argOuts_19_bits;
  assign regs_21_io_init = 64'h0;
  assign regs_21_io_enable = 1'h1;
  assign regs_21_clock = clock;
  assign regs_21_reset = reset;
  assign regs_22_io_in = io_argOuts_20_bits;
  assign regs_22_io_init = 64'h0;
  assign regs_22_io_enable = 1'h1;
  assign regs_22_clock = clock;
  assign regs_22_reset = reset;
  assign regs_23_io_in = io_argOuts_21_bits;
  assign regs_23_io_init = 64'h0;
  assign regs_23_io_enable = 1'h1;
  assign regs_23_clock = clock;
  assign regs_23_reset = reset;
  assign regs_24_io_in = io_argOuts_22_bits;
  assign regs_24_io_init = 64'h0;
  assign regs_24_io_enable = 1'h1;
  assign regs_24_clock = clock;
  assign regs_24_reset = reset;
  assign regs_25_io_in = io_argOuts_23_bits;
  assign regs_25_io_init = 64'h0;
  assign regs_25_io_enable = 1'h1;
  assign regs_25_clock = clock;
  assign regs_25_reset = reset;
  assign regs_26_io_in = io_argOuts_24_bits;
  assign regs_26_io_init = 64'h0;
  assign regs_26_io_enable = 1'h1;
  assign regs_26_clock = clock;
  assign regs_26_reset = reset;
  assign regs_27_io_in = io_argOuts_25_bits;
  assign regs_27_io_init = 64'h0;
  assign regs_27_io_enable = 1'h1;
  assign regs_27_clock = clock;
  assign regs_27_reset = reset;
  assign regs_28_io_in = io_argOuts_26_bits;
  assign regs_28_io_init = 64'h0;
  assign regs_28_io_enable = 1'h1;
  assign regs_28_clock = clock;
  assign regs_28_reset = reset;
  assign regs_29_io_in = io_argOuts_27_bits;
  assign regs_29_io_init = 64'h0;
  assign regs_29_io_enable = 1'h1;
  assign regs_29_clock = clock;
  assign regs_29_reset = reset;
  assign regs_30_io_in = io_argOuts_28_bits;
  assign regs_30_io_init = 64'h0;
  assign regs_30_io_enable = 1'h1;
  assign regs_30_clock = clock;
  assign regs_30_reset = reset;
  assign regs_31_io_in = io_argOuts_29_bits;
  assign regs_31_io_init = 64'h0;
  assign regs_31_io_enable = 1'h1;
  assign regs_31_clock = clock;
  assign regs_31_reset = reset;
  assign regs_32_io_in = io_argOuts_30_bits;
  assign regs_32_io_init = 64'h0;
  assign regs_32_io_enable = 1'h1;
  assign regs_32_clock = clock;
  assign regs_32_reset = reset;
  assign regs_33_io_in = io_argOuts_31_bits;
  assign regs_33_io_init = 64'h0;
  assign regs_33_io_enable = 1'h1;
  assign regs_33_clock = clock;
  assign regs_33_reset = reset;
  assign regs_34_io_in = io_argOuts_32_bits;
  assign regs_34_io_init = 64'h0;
  assign regs_34_io_enable = 1'h1;
  assign regs_34_clock = clock;
  assign regs_34_reset = reset;
  assign regs_35_io_in = io_argOuts_33_bits;
  assign regs_35_io_init = 64'h0;
  assign regs_35_io_enable = 1'h1;
  assign regs_35_clock = clock;
  assign regs_35_reset = reset;
  assign regs_36_io_in = io_argOuts_34_bits;
  assign regs_36_io_init = 64'h0;
  assign regs_36_io_enable = 1'h1;
  assign regs_36_clock = clock;
  assign regs_36_reset = reset;
  assign regs_37_io_in = io_argOuts_35_bits;
  assign regs_37_io_init = 64'h0;
  assign regs_37_io_enable = 1'h1;
  assign regs_37_clock = clock;
  assign regs_37_reset = reset;
  assign regs_38_io_in = io_argOuts_36_bits;
  assign regs_38_io_init = 64'h0;
  assign regs_38_io_enable = 1'h1;
  assign regs_38_clock = clock;
  assign regs_38_reset = reset;
  assign regs_39_io_in = io_argOuts_37_bits;
  assign regs_39_io_init = 64'h0;
  assign regs_39_io_enable = 1'h1;
  assign regs_39_clock = clock;
  assign regs_39_reset = reset;
  assign regs_40_io_in = io_argOuts_38_bits;
  assign regs_40_io_init = 64'h0;
  assign regs_40_io_enable = 1'h1;
  assign regs_40_clock = clock;
  assign regs_40_reset = reset;
  assign regs_41_io_in = io_argOuts_39_bits;
  assign regs_41_io_init = 64'h0;
  assign regs_41_io_enable = 1'h1;
  assign regs_41_clock = clock;
  assign regs_41_reset = reset;
  assign regs_42_io_in = io_argOuts_40_bits;
  assign regs_42_io_init = 64'h0;
  assign regs_42_io_enable = 1'h1;
  assign regs_42_clock = clock;
  assign regs_42_reset = reset;
  assign regs_43_io_in = io_argOuts_41_bits;
  assign regs_43_io_init = 64'h0;
  assign regs_43_io_enable = 1'h1;
  assign regs_43_clock = clock;
  assign regs_43_reset = reset;
  assign regs_44_io_in = io_argOuts_42_bits;
  assign regs_44_io_init = 64'h0;
  assign regs_44_io_enable = 1'h1;
  assign regs_44_clock = clock;
  assign regs_44_reset = reset;
  assign regs_45_io_in = io_argOuts_43_bits;
  assign regs_45_io_init = 64'h0;
  assign regs_45_io_enable = 1'h1;
  assign regs_45_clock = clock;
  assign regs_45_reset = reset;
  assign regs_46_io_in = io_argOuts_44_bits;
  assign regs_46_io_init = 64'h0;
  assign regs_46_io_enable = 1'h1;
  assign regs_46_clock = clock;
  assign regs_46_reset = reset;
  assign regs_47_io_in = io_argOuts_45_bits;
  assign regs_47_io_init = 64'h0;
  assign regs_47_io_enable = 1'h1;
  assign regs_47_clock = clock;
  assign regs_47_reset = reset;
  assign regs_48_io_in = io_argOuts_46_bits;
  assign regs_48_io_init = 64'h0;
  assign regs_48_io_enable = 1'h1;
  assign regs_48_clock = clock;
  assign regs_48_reset = reset;
  assign regs_49_io_in = io_argOuts_47_bits;
  assign regs_49_io_init = 64'h0;
  assign regs_49_io_enable = 1'h1;
  assign regs_49_clock = clock;
  assign regs_49_reset = reset;
  assign regs_50_io_in = io_argOuts_48_bits;
  assign regs_50_io_init = 64'h0;
  assign regs_50_io_enable = 1'h1;
  assign regs_50_clock = clock;
  assign regs_50_reset = reset;
  assign regs_51_io_in = io_argOuts_49_bits;
  assign regs_51_io_init = 64'h0;
  assign regs_51_io_enable = 1'h1;
  assign regs_51_clock = clock;
  assign regs_51_reset = reset;
  assign regs_52_io_in = io_argOuts_50_bits;
  assign regs_52_io_init = 64'h0;
  assign regs_52_io_enable = 1'h1;
  assign regs_52_clock = clock;
  assign regs_52_reset = reset;
  assign regs_53_io_in = io_argOuts_51_bits;
  assign regs_53_io_init = 64'h0;
  assign regs_53_io_enable = 1'h1;
  assign regs_53_clock = clock;
  assign regs_53_reset = reset;
  assign regs_54_io_in = io_argOuts_52_bits;
  assign regs_54_io_init = 64'h0;
  assign regs_54_io_enable = 1'h1;
  assign regs_54_clock = clock;
  assign regs_54_reset = reset;
  assign regs_55_io_in = io_argOuts_53_bits;
  assign regs_55_io_init = 64'h0;
  assign regs_55_io_enable = 1'h1;
  assign regs_55_clock = clock;
  assign regs_55_reset = reset;
  assign regs_56_io_in = io_argOuts_54_bits;
  assign regs_56_io_init = 64'h0;
  assign regs_56_io_enable = 1'h1;
  assign regs_56_clock = clock;
  assign regs_56_reset = reset;
  assign regs_57_io_in = io_argOuts_55_bits;
  assign regs_57_io_init = 64'h0;
  assign regs_57_io_enable = 1'h1;
  assign regs_57_clock = clock;
  assign regs_57_reset = reset;
  assign regs_58_io_in = io_argOuts_56_bits;
  assign regs_58_io_init = 64'h0;
  assign regs_58_io_enable = 1'h1;
  assign regs_58_clock = clock;
  assign regs_58_reset = reset;
  assign regs_59_io_in = io_argOuts_57_bits;
  assign regs_59_io_init = 64'h0;
  assign regs_59_io_enable = 1'h1;
  assign regs_59_clock = clock;
  assign regs_59_reset = reset;
  assign regs_60_io_in = io_argOuts_58_bits;
  assign regs_60_io_init = 64'h0;
  assign regs_60_io_enable = 1'h1;
  assign regs_60_clock = clock;
  assign regs_60_reset = reset;
  assign regs_61_io_in = io_argOuts_59_bits;
  assign regs_61_io_init = 64'h0;
  assign regs_61_io_enable = 1'h1;
  assign regs_61_clock = clock;
  assign regs_61_reset = reset;
  assign regs_62_io_in = io_argOuts_60_bits;
  assign regs_62_io_init = 64'h0;
  assign regs_62_io_enable = 1'h1;
  assign regs_62_clock = clock;
  assign regs_62_reset = reset;
  assign regs_63_io_in = 64'h0;
  assign regs_63_io_init = 64'h0;
  assign regs_63_io_enable = 1'h1;
  assign regs_63_clock = clock;
  assign regs_63_reset = reset;
  assign regs_64_io_in = 64'h0;
  assign regs_64_io_init = 64'h0;
  assign regs_64_io_enable = 1'h1;
  assign regs_64_clock = clock;
  assign regs_64_reset = reset;
  assign regs_65_io_in = 64'h0;
  assign regs_65_io_init = 64'h0;
  assign regs_65_io_enable = 1'h1;
  assign regs_65_clock = clock;
  assign regs_65_reset = reset;
  assign regs_66_io_in = 64'h0;
  assign regs_66_io_init = 64'h0;
  assign regs_66_io_enable = 1'h1;
  assign regs_66_clock = clock;
  assign regs_66_reset = reset;
  assign regs_67_io_in = 64'h0;
  assign regs_67_io_init = 64'h0;
  assign regs_67_io_enable = 1'h1;
  assign regs_67_clock = clock;
  assign regs_67_reset = reset;
  assign regs_68_io_in = 64'h0;
  assign regs_68_io_init = 64'h0;
  assign regs_68_io_enable = 1'h1;
  assign regs_68_clock = clock;
  assign regs_68_reset = reset;
  assign regs_69_io_in = 64'h0;
  assign regs_69_io_init = 64'h0;
  assign regs_69_io_enable = 1'h1;
  assign regs_69_clock = clock;
  assign regs_69_reset = reset;
  assign regs_70_io_in = 64'h0;
  assign regs_70_io_init = 64'h0;
  assign regs_70_io_enable = 1'h1;
  assign regs_70_clock = clock;
  assign regs_70_reset = reset;
  assign regs_71_io_in = 64'h0;
  assign regs_71_io_init = 64'h0;
  assign regs_71_io_enable = 1'h1;
  assign regs_71_clock = clock;
  assign regs_71_reset = reset;
  assign regs_72_io_in = 64'h0;
  assign regs_72_io_init = 64'h0;
  assign regs_72_io_enable = 1'h1;
  assign regs_72_clock = clock;
  assign regs_72_reset = reset;
  assign regs_73_io_in = 64'h0;
  assign regs_73_io_init = 64'h0;
  assign regs_73_io_enable = 1'h1;
  assign regs_73_clock = clock;
  assign regs_73_reset = reset;
  assign regs_74_io_in = 64'h0;
  assign regs_74_io_init = 64'h0;
  assign regs_74_io_enable = 1'h1;
  assign regs_74_clock = clock;
  assign regs_74_reset = reset;
  assign regs_75_io_in = 64'h0;
  assign regs_75_io_init = 64'h0;
  assign regs_75_io_enable = 1'h1;
  assign regs_75_clock = clock;
  assign regs_75_reset = reset;
  assign regs_76_io_in = 64'h0;
  assign regs_76_io_init = 64'h0;
  assign regs_76_io_enable = 1'h1;
  assign regs_76_clock = clock;
  assign regs_76_reset = reset;
  assign regs_77_io_in = 64'h0;
  assign regs_77_io_init = 64'h0;
  assign regs_77_io_enable = 1'h1;
  assign regs_77_clock = clock;
  assign regs_77_reset = reset;
  assign regs_78_io_in = 64'h0;
  assign regs_78_io_init = 64'h0;
  assign regs_78_io_enable = 1'h1;
  assign regs_78_clock = clock;
  assign regs_78_reset = reset;
  assign regs_79_io_in = 64'h0;
  assign regs_79_io_init = 64'h0;
  assign regs_79_io_enable = 1'h1;
  assign regs_79_clock = clock;
  assign regs_79_reset = reset;
  assign regs_80_io_in = 64'h0;
  assign regs_80_io_init = 64'h0;
  assign regs_80_io_enable = 1'h1;
  assign regs_80_clock = clock;
  assign regs_80_reset = reset;
  assign regs_81_io_in = 64'h0;
  assign regs_81_io_init = 64'h0;
  assign regs_81_io_enable = 1'h1;
  assign regs_81_clock = clock;
  assign regs_81_reset = reset;
  assign regs_82_io_in = 64'h0;
  assign regs_82_io_init = 64'h0;
  assign regs_82_io_enable = 1'h1;
  assign regs_82_clock = clock;
  assign regs_82_reset = reset;
  assign regs_83_io_in = 64'h0;
  assign regs_83_io_init = 64'h0;
  assign regs_83_io_enable = 1'h1;
  assign regs_83_clock = clock;
  assign regs_83_reset = reset;
  assign regs_84_io_in = 64'h0;
  assign regs_84_io_init = 64'h0;
  assign regs_84_io_enable = 1'h1;
  assign regs_84_clock = clock;
  assign regs_84_reset = reset;
  assign regs_85_io_in = 64'h0;
  assign regs_85_io_init = 64'h0;
  assign regs_85_io_enable = 1'h1;
  assign regs_85_clock = clock;
  assign regs_85_reset = reset;
  assign regs_86_io_in = 64'h0;
  assign regs_86_io_init = 64'h0;
  assign regs_86_io_enable = 1'h1;
  assign regs_86_clock = clock;
  assign regs_86_reset = reset;
  assign regs_87_io_in = 64'h0;
  assign regs_87_io_init = 64'h0;
  assign regs_87_io_enable = 1'h1;
  assign regs_87_clock = clock;
  assign regs_87_reset = reset;
  assign regs_88_io_in = 64'h0;
  assign regs_88_io_init = 64'h0;
  assign regs_88_io_enable = 1'h1;
  assign regs_88_clock = clock;
  assign regs_88_reset = reset;
  assign regs_89_io_in = 64'h0;
  assign regs_89_io_init = 64'h0;
  assign regs_89_io_enable = 1'h1;
  assign regs_89_clock = clock;
  assign regs_89_reset = reset;
  assign regs_90_io_in = 64'h0;
  assign regs_90_io_init = 64'h0;
  assign regs_90_io_enable = 1'h1;
  assign regs_90_clock = clock;
  assign regs_90_reset = reset;
  assign regs_91_io_in = 64'h0;
  assign regs_91_io_init = 64'h0;
  assign regs_91_io_enable = 1'h1;
  assign regs_91_clock = clock;
  assign regs_91_reset = reset;
  assign regs_92_io_in = 64'h0;
  assign regs_92_io_init = 64'h0;
  assign regs_92_io_enable = 1'h1;
  assign regs_92_clock = clock;
  assign regs_92_reset = reset;
  assign regs_93_io_in = 64'h0;
  assign regs_93_io_init = 64'h0;
  assign regs_93_io_enable = 1'h1;
  assign regs_93_clock = clock;
  assign regs_93_reset = reset;
  assign regs_94_io_in = 64'h0;
  assign regs_94_io_init = 64'h0;
  assign regs_94_io_enable = 1'h1;
  assign regs_94_clock = clock;
  assign regs_94_reset = reset;
  assign regs_95_io_in = 64'h0;
  assign regs_95_io_init = 64'h0;
  assign regs_95_io_enable = 1'h1;
  assign regs_95_clock = clock;
  assign regs_95_reset = reset;
  assign regs_96_io_in = 64'h0;
  assign regs_96_io_init = 64'h0;
  assign regs_96_io_enable = 1'h1;
  assign regs_96_clock = clock;
  assign regs_96_reset = reset;
  assign regs_97_io_in = 64'h0;
  assign regs_97_io_init = 64'h0;
  assign regs_97_io_enable = 1'h1;
  assign regs_97_clock = clock;
  assign regs_97_reset = reset;
  assign regs_98_io_in = 64'h0;
  assign regs_98_io_init = 64'h0;
  assign regs_98_io_enable = 1'h1;
  assign regs_98_clock = clock;
  assign regs_98_reset = reset;
  assign regs_99_io_in = 64'h0;
  assign regs_99_io_init = 64'h0;
  assign regs_99_io_enable = 1'h1;
  assign regs_99_clock = clock;
  assign regs_99_reset = reset;
  assign regs_100_io_in = 64'h0;
  assign regs_100_io_init = 64'h0;
  assign regs_100_io_enable = 1'h1;
  assign regs_100_clock = clock;
  assign regs_100_reset = reset;
  assign regs_101_io_in = 64'h0;
  assign regs_101_io_init = 64'h0;
  assign regs_101_io_enable = 1'h1;
  assign regs_101_clock = clock;
  assign regs_101_reset = reset;
  assign regs_102_io_in = 64'h0;
  assign regs_102_io_init = 64'h0;
  assign regs_102_io_enable = 1'h1;
  assign regs_102_clock = clock;
  assign regs_102_reset = reset;
  assign regs_103_io_in = 64'h0;
  assign regs_103_io_init = 64'h0;
  assign regs_103_io_enable = 1'h1;
  assign regs_103_clock = clock;
  assign regs_103_reset = reset;
  assign regs_104_io_in = 64'h0;
  assign regs_104_io_init = 64'h0;
  assign regs_104_io_enable = 1'h1;
  assign regs_104_clock = clock;
  assign regs_104_reset = reset;
  assign regs_105_io_in = 64'h0;
  assign regs_105_io_init = 64'h0;
  assign regs_105_io_enable = 1'h1;
  assign regs_105_clock = clock;
  assign regs_105_reset = reset;
  assign regs_106_io_in = 64'h0;
  assign regs_106_io_init = 64'h0;
  assign regs_106_io_enable = 1'h1;
  assign regs_106_clock = clock;
  assign regs_106_reset = reset;
  assign regs_107_io_in = 64'h0;
  assign regs_107_io_init = 64'h0;
  assign regs_107_io_enable = 1'h1;
  assign regs_107_clock = clock;
  assign regs_107_reset = reset;
  assign regs_108_io_in = 64'h0;
  assign regs_108_io_init = 64'h0;
  assign regs_108_io_enable = 1'h1;
  assign regs_108_clock = clock;
  assign regs_108_reset = reset;
  assign regs_109_io_in = 64'h0;
  assign regs_109_io_init = 64'h0;
  assign regs_109_io_enable = 1'h1;
  assign regs_109_clock = clock;
  assign regs_109_reset = reset;
  assign regs_110_io_in = 64'h0;
  assign regs_110_io_init = 64'h0;
  assign regs_110_io_enable = 1'h1;
  assign regs_110_clock = clock;
  assign regs_110_reset = reset;
  assign regs_111_io_in = 64'h0;
  assign regs_111_io_init = 64'h0;
  assign regs_111_io_enable = 1'h1;
  assign regs_111_clock = clock;
  assign regs_111_reset = reset;
  assign regs_112_io_in = 64'h0;
  assign regs_112_io_init = 64'h0;
  assign regs_112_io_enable = 1'h1;
  assign regs_112_clock = clock;
  assign regs_112_reset = reset;
  assign regs_113_io_in = 64'h0;
  assign regs_113_io_init = 64'h0;
  assign regs_113_io_enable = 1'h1;
  assign regs_113_clock = clock;
  assign regs_113_reset = reset;
  assign regs_114_io_in = 64'h0;
  assign regs_114_io_init = 64'h0;
  assign regs_114_io_enable = 1'h1;
  assign regs_114_clock = clock;
  assign regs_114_reset = reset;
  assign regs_115_io_in = 64'h0;
  assign regs_115_io_init = 64'h0;
  assign regs_115_io_enable = 1'h1;
  assign regs_115_clock = clock;
  assign regs_115_reset = reset;
  assign regs_116_io_in = 64'h0;
  assign regs_116_io_init = 64'h0;
  assign regs_116_io_enable = 1'h1;
  assign regs_116_clock = clock;
  assign regs_116_reset = reset;
  assign regs_117_io_in = 64'h0;
  assign regs_117_io_init = 64'h0;
  assign regs_117_io_enable = 1'h1;
  assign regs_117_clock = clock;
  assign regs_117_reset = reset;
  assign regs_118_io_in = 64'h0;
  assign regs_118_io_init = 64'h0;
  assign regs_118_io_enable = 1'h1;
  assign regs_118_clock = clock;
  assign regs_118_reset = reset;
  assign regs_119_io_in = 64'h0;
  assign regs_119_io_init = 64'h0;
  assign regs_119_io_enable = 1'h1;
  assign regs_119_clock = clock;
  assign regs_119_reset = reset;
  assign regs_120_io_in = 64'h0;
  assign regs_120_io_init = 64'h0;
  assign regs_120_io_enable = 1'h1;
  assign regs_120_clock = clock;
  assign regs_120_reset = reset;
  assign regs_121_io_in = 64'h0;
  assign regs_121_io_init = 64'h0;
  assign regs_121_io_enable = 1'h1;
  assign regs_121_clock = clock;
  assign regs_121_reset = reset;
  assign regs_122_io_in = 64'h0;
  assign regs_122_io_init = 64'h0;
  assign regs_122_io_enable = 1'h1;
  assign regs_122_clock = clock;
  assign regs_122_reset = reset;
  assign regs_123_io_in = 64'h0;
  assign regs_123_io_init = 64'h0;
  assign regs_123_io_enable = 1'h1;
  assign regs_123_clock = clock;
  assign regs_123_reset = reset;
  assign regs_124_io_in = 64'h0;
  assign regs_124_io_init = 64'h0;
  assign regs_124_io_enable = 1'h1;
  assign regs_124_clock = clock;
  assign regs_124_reset = reset;
  assign regs_125_io_in = 64'h0;
  assign regs_125_io_init = 64'h0;
  assign regs_125_io_enable = 1'h1;
  assign regs_125_clock = clock;
  assign regs_125_reset = reset;
  assign regs_126_io_in = 64'h0;
  assign regs_126_io_init = 64'h0;
  assign regs_126_io_enable = 1'h1;
  assign regs_126_clock = clock;
  assign regs_126_reset = reset;
  assign regs_127_io_in = 64'h0;
  assign regs_127_io_init = 64'h0;
  assign regs_127_io_enable = 1'h1;
  assign regs_127_clock = clock;
  assign regs_127_reset = reset;
  assign regs_128_io_in = 64'h0;
  assign regs_128_io_init = 64'h0;
  assign regs_128_io_enable = 1'h1;
  assign regs_128_clock = clock;
  assign regs_128_reset = reset;
  assign regs_129_io_in = 64'h0;
  assign regs_129_io_init = 64'h0;
  assign regs_129_io_enable = 1'h1;
  assign regs_129_clock = clock;
  assign regs_129_reset = reset;
  assign regs_130_io_in = 64'h0;
  assign regs_130_io_init = 64'h0;
  assign regs_130_io_enable = 1'h1;
  assign regs_130_clock = clock;
  assign regs_130_reset = reset;
  assign regs_131_io_in = 64'h0;
  assign regs_131_io_init = 64'h0;
  assign regs_131_io_enable = 1'h1;
  assign regs_131_clock = clock;
  assign regs_131_reset = reset;
  assign regs_132_io_in = 64'h0;
  assign regs_132_io_init = 64'h0;
  assign regs_132_io_enable = 1'h1;
  assign regs_132_clock = clock;
  assign regs_132_reset = reset;
  assign regs_133_io_in = 64'h0;
  assign regs_133_io_init = 64'h0;
  assign regs_133_io_enable = 1'h1;
  assign regs_133_clock = clock;
  assign regs_133_reset = reset;
  assign regs_134_io_in = 64'h0;
  assign regs_134_io_init = 64'h0;
  assign regs_134_io_enable = 1'h1;
  assign regs_134_clock = clock;
  assign regs_134_reset = reset;
  assign regs_135_io_in = 64'h0;
  assign regs_135_io_init = 64'h0;
  assign regs_135_io_enable = 1'h1;
  assign regs_135_clock = clock;
  assign regs_135_reset = reset;
  assign regs_136_io_in = 64'h0;
  assign regs_136_io_init = 64'h0;
  assign regs_136_io_enable = 1'h1;
  assign regs_136_clock = clock;
  assign regs_136_reset = reset;
  assign regs_137_io_in = 64'h0;
  assign regs_137_io_init = 64'h0;
  assign regs_137_io_enable = 1'h1;
  assign regs_137_clock = clock;
  assign regs_137_reset = reset;
  assign regs_138_io_in = 64'h0;
  assign regs_138_io_init = 64'h0;
  assign regs_138_io_enable = 1'h1;
  assign regs_138_clock = clock;
  assign regs_138_reset = reset;
  assign regs_139_io_in = 64'h0;
  assign regs_139_io_init = 64'h0;
  assign regs_139_io_enable = 1'h1;
  assign regs_139_clock = clock;
  assign regs_139_reset = reset;
  assign regs_140_io_in = 64'h0;
  assign regs_140_io_init = 64'h0;
  assign regs_140_io_enable = 1'h1;
  assign regs_140_clock = clock;
  assign regs_140_reset = reset;
  assign regs_141_io_in = 64'h0;
  assign regs_141_io_init = 64'h0;
  assign regs_141_io_enable = 1'h1;
  assign regs_141_clock = clock;
  assign regs_141_reset = reset;
  assign regs_142_io_in = 64'h0;
  assign regs_142_io_init = 64'h0;
  assign regs_142_io_enable = 1'h1;
  assign regs_142_clock = clock;
  assign regs_142_reset = reset;
  assign regs_143_io_in = 64'h0;
  assign regs_143_io_init = 64'h0;
  assign regs_143_io_enable = 1'h1;
  assign regs_143_clock = clock;
  assign regs_143_reset = reset;
  assign regs_144_io_in = 64'h0;
  assign regs_144_io_init = 64'h0;
  assign regs_144_io_enable = 1'h1;
  assign regs_144_clock = clock;
  assign regs_144_reset = reset;
  assign regs_145_io_in = 64'h0;
  assign regs_145_io_init = 64'h0;
  assign regs_145_io_enable = 1'h1;
  assign regs_145_clock = clock;
  assign regs_145_reset = reset;
  assign regs_146_io_in = 64'h0;
  assign regs_146_io_init = 64'h0;
  assign regs_146_io_enable = 1'h1;
  assign regs_146_clock = clock;
  assign regs_146_reset = reset;
  assign regs_147_io_in = 64'h0;
  assign regs_147_io_init = 64'h0;
  assign regs_147_io_enable = 1'h1;
  assign regs_147_clock = clock;
  assign regs_147_reset = reset;
  assign regs_148_io_in = 64'h0;
  assign regs_148_io_init = 64'h0;
  assign regs_148_io_enable = 1'h1;
  assign regs_148_clock = clock;
  assign regs_148_reset = reset;
  assign regs_149_io_in = 64'h0;
  assign regs_149_io_init = 64'h0;
  assign regs_149_io_enable = 1'h1;
  assign regs_149_clock = clock;
  assign regs_149_reset = reset;
  assign regs_150_io_in = 64'h0;
  assign regs_150_io_init = 64'h0;
  assign regs_150_io_enable = 1'h1;
  assign regs_150_clock = clock;
  assign regs_150_reset = reset;
  assign regs_151_io_in = 64'h0;
  assign regs_151_io_init = 64'h0;
  assign regs_151_io_enable = 1'h1;
  assign regs_151_clock = clock;
  assign regs_151_reset = reset;
  assign regs_152_io_in = 64'h0;
  assign regs_152_io_init = 64'h0;
  assign regs_152_io_enable = 1'h1;
  assign regs_152_clock = clock;
  assign regs_152_reset = reset;
  assign regs_153_io_in = 64'h0;
  assign regs_153_io_init = 64'h0;
  assign regs_153_io_enable = 1'h1;
  assign regs_153_clock = clock;
  assign regs_153_reset = reset;
  assign regs_154_io_in = 64'h0;
  assign regs_154_io_init = 64'h0;
  assign regs_154_io_enable = 1'h1;
  assign regs_154_clock = clock;
  assign regs_154_reset = reset;
  assign regs_155_io_in = 64'h0;
  assign regs_155_io_init = 64'h0;
  assign regs_155_io_enable = 1'h1;
  assign regs_155_clock = clock;
  assign regs_155_reset = reset;
  assign regs_156_io_in = 64'h0;
  assign regs_156_io_init = 64'h0;
  assign regs_156_io_enable = 1'h1;
  assign regs_156_clock = clock;
  assign regs_156_reset = reset;
  assign regs_157_io_in = 64'h0;
  assign regs_157_io_init = 64'h0;
  assign regs_157_io_enable = 1'h1;
  assign regs_157_clock = clock;
  assign regs_157_reset = reset;
  assign regs_158_io_in = 64'h0;
  assign regs_158_io_init = 64'h0;
  assign regs_158_io_enable = 1'h1;
  assign regs_158_clock = clock;
  assign regs_158_reset = reset;
  assign regs_159_io_in = 64'h0;
  assign regs_159_io_init = 64'h0;
  assign regs_159_io_enable = 1'h1;
  assign regs_159_clock = clock;
  assign regs_159_reset = reset;
  assign regs_160_io_in = 64'h0;
  assign regs_160_io_init = 64'h0;
  assign regs_160_io_enable = 1'h1;
  assign regs_160_clock = clock;
  assign regs_160_reset = reset;
  assign regs_161_io_in = 64'h0;
  assign regs_161_io_init = 64'h0;
  assign regs_161_io_enable = 1'h1;
  assign regs_161_clock = clock;
  assign regs_161_reset = reset;
  assign regs_162_io_in = 64'h0;
  assign regs_162_io_init = 64'h0;
  assign regs_162_io_enable = 1'h1;
  assign regs_162_clock = clock;
  assign regs_162_reset = reset;
  assign regs_163_io_in = 64'h0;
  assign regs_163_io_init = 64'h0;
  assign regs_163_io_enable = 1'h1;
  assign regs_163_clock = clock;
  assign regs_163_reset = reset;
  assign regs_164_io_in = 64'h0;
  assign regs_164_io_init = 64'h0;
  assign regs_164_io_enable = 1'h1;
  assign regs_164_clock = clock;
  assign regs_164_reset = reset;
  assign regs_165_io_in = 64'h0;
  assign regs_165_io_init = 64'h0;
  assign regs_165_io_enable = 1'h1;
  assign regs_165_clock = clock;
  assign regs_165_reset = reset;
  assign regs_166_io_in = 64'h0;
  assign regs_166_io_init = 64'h0;
  assign regs_166_io_enable = 1'h1;
  assign regs_166_clock = clock;
  assign regs_166_reset = reset;
  assign regs_167_io_in = 64'h0;
  assign regs_167_io_init = 64'h0;
  assign regs_167_io_enable = 1'h1;
  assign regs_167_clock = clock;
  assign regs_167_reset = reset;
  assign regs_168_io_in = 64'h0;
  assign regs_168_io_init = 64'h0;
  assign regs_168_io_enable = 1'h1;
  assign regs_168_clock = clock;
  assign regs_168_reset = reset;
  assign regs_169_io_in = 64'h0;
  assign regs_169_io_init = 64'h0;
  assign regs_169_io_enable = 1'h1;
  assign regs_169_clock = clock;
  assign regs_169_reset = reset;
  assign regs_170_io_in = 64'h0;
  assign regs_170_io_init = 64'h0;
  assign regs_170_io_enable = 1'h1;
  assign regs_170_clock = clock;
  assign regs_170_reset = reset;
  assign regs_171_io_in = 64'h0;
  assign regs_171_io_init = 64'h0;
  assign regs_171_io_enable = 1'h1;
  assign regs_171_clock = clock;
  assign regs_171_reset = reset;
  assign regs_172_io_in = 64'h0;
  assign regs_172_io_init = 64'h0;
  assign regs_172_io_enable = 1'h1;
  assign regs_172_clock = clock;
  assign regs_172_reset = reset;
  assign regs_173_io_in = 64'h0;
  assign regs_173_io_init = 64'h0;
  assign regs_173_io_enable = 1'h1;
  assign regs_173_clock = clock;
  assign regs_173_reset = reset;
  assign regs_174_io_in = 64'h0;
  assign regs_174_io_init = 64'h0;
  assign regs_174_io_enable = 1'h1;
  assign regs_174_clock = clock;
  assign regs_174_reset = reset;
  assign regs_175_io_in = 64'h0;
  assign regs_175_io_init = 64'h0;
  assign regs_175_io_enable = 1'h1;
  assign regs_175_clock = clock;
  assign regs_175_reset = reset;
  assign regs_176_io_in = 64'h0;
  assign regs_176_io_init = 64'h0;
  assign regs_176_io_enable = 1'h1;
  assign regs_176_clock = clock;
  assign regs_176_reset = reset;
  assign regs_177_io_in = 64'h0;
  assign regs_177_io_init = 64'h0;
  assign regs_177_io_enable = 1'h1;
  assign regs_177_clock = clock;
  assign regs_177_reset = reset;
  assign regs_178_io_in = 64'h0;
  assign regs_178_io_init = 64'h0;
  assign regs_178_io_enable = 1'h1;
  assign regs_178_clock = clock;
  assign regs_178_reset = reset;
  assign regs_179_io_in = 64'h0;
  assign regs_179_io_init = 64'h0;
  assign regs_179_io_enable = 1'h1;
  assign regs_179_clock = clock;
  assign regs_179_reset = reset;
  assign regs_180_io_in = 64'h0;
  assign regs_180_io_init = 64'h0;
  assign regs_180_io_enable = 1'h1;
  assign regs_180_clock = clock;
  assign regs_180_reset = reset;
  assign regs_181_io_in = 64'h0;
  assign regs_181_io_init = 64'h0;
  assign regs_181_io_enable = 1'h1;
  assign regs_181_clock = clock;
  assign regs_181_reset = reset;
  assign regs_182_io_in = 64'h0;
  assign regs_182_io_init = 64'h0;
  assign regs_182_io_enable = 1'h1;
  assign regs_182_clock = clock;
  assign regs_182_reset = reset;
  assign regs_183_io_in = 64'h0;
  assign regs_183_io_init = 64'h0;
  assign regs_183_io_enable = 1'h1;
  assign regs_183_clock = clock;
  assign regs_183_reset = reset;
  assign regs_184_io_in = 64'h0;
  assign regs_184_io_init = 64'h0;
  assign regs_184_io_enable = 1'h1;
  assign regs_184_clock = clock;
  assign regs_184_reset = reset;
  assign regs_185_io_in = 64'h0;
  assign regs_185_io_init = 64'h0;
  assign regs_185_io_enable = 1'h1;
  assign regs_185_clock = clock;
  assign regs_185_reset = reset;
  assign regs_186_io_in = 64'h0;
  assign regs_186_io_init = 64'h0;
  assign regs_186_io_enable = 1'h1;
  assign regs_186_clock = clock;
  assign regs_186_reset = reset;
  assign regs_187_io_in = 64'h0;
  assign regs_187_io_init = 64'h0;
  assign regs_187_io_enable = 1'h1;
  assign regs_187_clock = clock;
  assign regs_187_reset = reset;
  assign regs_188_io_in = 64'h0;
  assign regs_188_io_init = 64'h0;
  assign regs_188_io_enable = 1'h1;
  assign regs_188_clock = clock;
  assign regs_188_reset = reset;
  assign regs_189_io_in = 64'h0;
  assign regs_189_io_init = 64'h0;
  assign regs_189_io_enable = 1'h1;
  assign regs_189_clock = clock;
  assign regs_189_reset = reset;
  assign regs_190_io_in = 64'h0;
  assign regs_190_io_init = 64'h0;
  assign regs_190_io_enable = 1'h1;
  assign regs_190_clock = clock;
  assign regs_190_reset = reset;
  assign regs_191_io_in = 64'h0;
  assign regs_191_io_init = 64'h0;
  assign regs_191_io_enable = 1'h1;
  assign regs_191_clock = clock;
  assign regs_191_reset = reset;
  assign regs_192_io_in = 64'h0;
  assign regs_192_io_init = 64'h0;
  assign regs_192_io_enable = 1'h1;
  assign regs_192_clock = clock;
  assign regs_192_reset = reset;
  assign regs_193_io_in = 64'h0;
  assign regs_193_io_init = 64'h0;
  assign regs_193_io_enable = 1'h1;
  assign regs_193_clock = clock;
  assign regs_193_reset = reset;
  assign regs_194_io_in = 64'h0;
  assign regs_194_io_init = 64'h0;
  assign regs_194_io_enable = 1'h1;
  assign regs_194_clock = clock;
  assign regs_194_reset = reset;
  assign regs_195_io_in = 64'h0;
  assign regs_195_io_init = 64'h0;
  assign regs_195_io_enable = 1'h1;
  assign regs_195_clock = clock;
  assign regs_195_reset = reset;
  assign regs_196_io_in = 64'h0;
  assign regs_196_io_init = 64'h0;
  assign regs_196_io_enable = 1'h1;
  assign regs_196_clock = clock;
  assign regs_196_reset = reset;
  assign regs_197_io_in = 64'h0;
  assign regs_197_io_init = 64'h0;
  assign regs_197_io_enable = 1'h1;
  assign regs_197_clock = clock;
  assign regs_197_reset = reset;
  assign regs_198_io_in = 64'h0;
  assign regs_198_io_init = 64'h0;
  assign regs_198_io_enable = 1'h1;
  assign regs_198_clock = clock;
  assign regs_198_reset = reset;
  assign regs_199_io_in = 64'h0;
  assign regs_199_io_init = 64'h0;
  assign regs_199_io_enable = 1'h1;
  assign regs_199_clock = clock;
  assign regs_199_reset = reset;
  assign regs_200_io_in = 64'h0;
  assign regs_200_io_init = 64'h0;
  assign regs_200_io_enable = 1'h1;
  assign regs_200_clock = clock;
  assign regs_200_reset = reset;
  assign regs_201_io_in = 64'h0;
  assign regs_201_io_init = 64'h0;
  assign regs_201_io_enable = 1'h1;
  assign regs_201_clock = clock;
  assign regs_201_reset = reset;
  assign regs_202_io_in = 64'h0;
  assign regs_202_io_init = 64'h0;
  assign regs_202_io_enable = 1'h1;
  assign regs_202_clock = clock;
  assign regs_202_reset = reset;
  assign regs_203_io_in = 64'h0;
  assign regs_203_io_init = 64'h0;
  assign regs_203_io_enable = 1'h1;
  assign regs_203_clock = clock;
  assign regs_203_reset = reset;
  assign regs_204_io_in = 64'h0;
  assign regs_204_io_init = 64'h0;
  assign regs_204_io_enable = 1'h1;
  assign regs_204_clock = clock;
  assign regs_204_reset = reset;
  assign regs_205_io_in = 64'h0;
  assign regs_205_io_init = 64'h0;
  assign regs_205_io_enable = 1'h1;
  assign regs_205_clock = clock;
  assign regs_205_reset = reset;
  assign regs_206_io_in = 64'h0;
  assign regs_206_io_init = 64'h0;
  assign regs_206_io_enable = 1'h1;
  assign regs_206_clock = clock;
  assign regs_206_reset = reset;
  assign regs_207_io_in = 64'h0;
  assign regs_207_io_init = 64'h0;
  assign regs_207_io_enable = 1'h1;
  assign regs_207_clock = clock;
  assign regs_207_reset = reset;
  assign regs_208_io_in = 64'h0;
  assign regs_208_io_init = 64'h0;
  assign regs_208_io_enable = 1'h1;
  assign regs_208_clock = clock;
  assign regs_208_reset = reset;
  assign regs_209_io_in = 64'h0;
  assign regs_209_io_init = 64'h0;
  assign regs_209_io_enable = 1'h1;
  assign regs_209_clock = clock;
  assign regs_209_reset = reset;
  assign regs_210_io_in = 64'h0;
  assign regs_210_io_init = 64'h0;
  assign regs_210_io_enable = 1'h1;
  assign regs_210_clock = clock;
  assign regs_210_reset = reset;
  assign regs_211_io_in = 64'h0;
  assign regs_211_io_init = 64'h0;
  assign regs_211_io_enable = 1'h1;
  assign regs_211_clock = clock;
  assign regs_211_reset = reset;
  assign regs_212_io_in = 64'h0;
  assign regs_212_io_init = 64'h0;
  assign regs_212_io_enable = 1'h1;
  assign regs_212_clock = clock;
  assign regs_212_reset = reset;
  assign regs_213_io_in = 64'h0;
  assign regs_213_io_init = 64'h0;
  assign regs_213_io_enable = 1'h1;
  assign regs_213_clock = clock;
  assign regs_213_reset = reset;
  assign regs_214_io_in = 64'h0;
  assign regs_214_io_init = 64'h0;
  assign regs_214_io_enable = 1'h1;
  assign regs_214_clock = clock;
  assign regs_214_reset = reset;
  assign regs_215_io_in = 64'h0;
  assign regs_215_io_init = 64'h0;
  assign regs_215_io_enable = 1'h1;
  assign regs_215_clock = clock;
  assign regs_215_reset = reset;
  assign regs_216_io_in = 64'h0;
  assign regs_216_io_init = 64'h0;
  assign regs_216_io_enable = 1'h1;
  assign regs_216_clock = clock;
  assign regs_216_reset = reset;
  assign regs_217_io_in = 64'h0;
  assign regs_217_io_init = 64'h0;
  assign regs_217_io_enable = 1'h1;
  assign regs_217_clock = clock;
  assign regs_217_reset = reset;
  assign regs_218_io_in = 64'h0;
  assign regs_218_io_init = 64'h0;
  assign regs_218_io_enable = 1'h1;
  assign regs_218_clock = clock;
  assign regs_218_reset = reset;
  assign regs_219_io_in = 64'h0;
  assign regs_219_io_init = 64'h0;
  assign regs_219_io_enable = 1'h1;
  assign regs_219_clock = clock;
  assign regs_219_reset = reset;
  assign regs_220_io_in = 64'h0;
  assign regs_220_io_init = 64'h0;
  assign regs_220_io_enable = 1'h1;
  assign regs_220_clock = clock;
  assign regs_220_reset = reset;
  assign regs_221_io_in = 64'h0;
  assign regs_221_io_init = 64'h0;
  assign regs_221_io_enable = 1'h1;
  assign regs_221_clock = clock;
  assign regs_221_reset = reset;
  assign regs_222_io_in = 64'h0;
  assign regs_222_io_init = 64'h0;
  assign regs_222_io_enable = 1'h1;
  assign regs_222_clock = clock;
  assign regs_222_reset = reset;
  assign regs_223_io_in = 64'h0;
  assign regs_223_io_init = 64'h0;
  assign regs_223_io_enable = 1'h1;
  assign regs_223_clock = clock;
  assign regs_223_reset = reset;
  assign regs_224_io_in = 64'h0;
  assign regs_224_io_init = 64'h0;
  assign regs_224_io_enable = 1'h1;
  assign regs_224_clock = clock;
  assign regs_224_reset = reset;
  assign regs_225_io_in = 64'h0;
  assign regs_225_io_init = 64'h0;
  assign regs_225_io_enable = 1'h1;
  assign regs_225_clock = clock;
  assign regs_225_reset = reset;
  assign regs_226_io_in = 64'h0;
  assign regs_226_io_init = 64'h0;
  assign regs_226_io_enable = 1'h1;
  assign regs_226_clock = clock;
  assign regs_226_reset = reset;
  assign regs_227_io_in = 64'h0;
  assign regs_227_io_init = 64'h0;
  assign regs_227_io_enable = 1'h1;
  assign regs_227_clock = clock;
  assign regs_227_reset = reset;
  assign regs_228_io_in = 64'h0;
  assign regs_228_io_init = 64'h0;
  assign regs_228_io_enable = 1'h1;
  assign regs_228_clock = clock;
  assign regs_228_reset = reset;
  assign regs_229_io_in = 64'h0;
  assign regs_229_io_init = 64'h0;
  assign regs_229_io_enable = 1'h1;
  assign regs_229_clock = clock;
  assign regs_229_reset = reset;
  assign regs_230_io_in = 64'h0;
  assign regs_230_io_init = 64'h0;
  assign regs_230_io_enable = 1'h1;
  assign regs_230_clock = clock;
  assign regs_230_reset = reset;
  assign regs_231_io_in = 64'h0;
  assign regs_231_io_init = 64'h0;
  assign regs_231_io_enable = 1'h1;
  assign regs_231_clock = clock;
  assign regs_231_reset = reset;
  assign regs_232_io_in = 64'h0;
  assign regs_232_io_init = 64'h0;
  assign regs_232_io_enable = 1'h1;
  assign regs_232_clock = clock;
  assign regs_232_reset = reset;
  assign regs_233_io_in = 64'h0;
  assign regs_233_io_init = 64'h0;
  assign regs_233_io_enable = 1'h1;
  assign regs_233_clock = clock;
  assign regs_233_reset = reset;
  assign regs_234_io_in = 64'h0;
  assign regs_234_io_init = 64'h0;
  assign regs_234_io_enable = 1'h1;
  assign regs_234_clock = clock;
  assign regs_234_reset = reset;
  assign regs_235_io_in = 64'h0;
  assign regs_235_io_init = 64'h0;
  assign regs_235_io_enable = 1'h1;
  assign regs_235_clock = clock;
  assign regs_235_reset = reset;
  assign rport_io_ins_0 = regOuts_0;
  assign rport_io_ins_1 = regOuts_1;
  assign rport_io_ins_2 = regOuts_2;
  assign rport_io_ins_3 = regOuts_3;
  assign rport_io_ins_4 = regOuts_4;
  assign rport_io_ins_5 = regOuts_5;
  assign rport_io_ins_6 = regOuts_6;
  assign rport_io_ins_7 = regOuts_7;
  assign rport_io_ins_8 = regOuts_8;
  assign rport_io_ins_9 = regOuts_9;
  assign rport_io_ins_10 = regOuts_10;
  assign rport_io_ins_11 = regOuts_11;
  assign rport_io_ins_12 = regOuts_12;
  assign rport_io_ins_13 = regOuts_13;
  assign rport_io_ins_14 = regOuts_14;
  assign rport_io_ins_15 = regOuts_15;
  assign rport_io_ins_16 = regOuts_16;
  assign rport_io_ins_17 = regOuts_17;
  assign rport_io_ins_18 = regOuts_18;
  assign rport_io_ins_19 = regOuts_19;
  assign rport_io_ins_20 = regOuts_20;
  assign rport_io_ins_21 = regOuts_21;
  assign rport_io_ins_22 = regOuts_22;
  assign rport_io_ins_23 = regOuts_23;
  assign rport_io_ins_24 = regOuts_24;
  assign rport_io_ins_25 = regOuts_25;
  assign rport_io_ins_26 = regOuts_26;
  assign rport_io_ins_27 = regOuts_27;
  assign rport_io_ins_28 = regOuts_28;
  assign rport_io_ins_29 = regOuts_29;
  assign rport_io_ins_30 = regOuts_30;
  assign rport_io_ins_31 = regOuts_31;
  assign rport_io_ins_32 = regOuts_32;
  assign rport_io_ins_33 = regOuts_33;
  assign rport_io_ins_34 = regOuts_34;
  assign rport_io_ins_35 = regOuts_35;
  assign rport_io_ins_36 = regOuts_36;
  assign rport_io_ins_37 = regOuts_37;
  assign rport_io_ins_38 = regOuts_38;
  assign rport_io_ins_39 = regOuts_39;
  assign rport_io_ins_40 = regOuts_40;
  assign rport_io_ins_41 = regOuts_41;
  assign rport_io_ins_42 = regOuts_42;
  assign rport_io_ins_43 = regOuts_43;
  assign rport_io_ins_44 = regOuts_44;
  assign rport_io_ins_45 = regOuts_45;
  assign rport_io_ins_46 = regOuts_46;
  assign rport_io_ins_47 = regOuts_47;
  assign rport_io_ins_48 = regOuts_48;
  assign rport_io_ins_49 = regOuts_49;
  assign rport_io_ins_50 = regOuts_50;
  assign rport_io_ins_51 = regOuts_51;
  assign rport_io_ins_52 = regOuts_52;
  assign rport_io_ins_53 = regOuts_53;
  assign rport_io_ins_54 = regOuts_54;
  assign rport_io_ins_55 = regOuts_55;
  assign rport_io_ins_56 = regOuts_56;
  assign rport_io_ins_57 = regOuts_57;
  assign rport_io_ins_58 = regOuts_58;
  assign rport_io_ins_59 = regOuts_59;
  assign rport_io_ins_60 = regOuts_60;
  assign rport_io_ins_61 = regOuts_61;
  assign rport_io_ins_62 = regOuts_62;
  assign rport_io_ins_63 = regOuts_63;
  assign rport_io_ins_64 = regOuts_64;
  assign rport_io_ins_65 = regOuts_65;
  assign rport_io_ins_66 = regOuts_66;
  assign rport_io_ins_67 = regOuts_67;
  assign rport_io_ins_68 = regOuts_68;
  assign rport_io_ins_69 = regOuts_69;
  assign rport_io_ins_70 = regOuts_70;
  assign rport_io_ins_71 = regOuts_71;
  assign rport_io_ins_72 = regOuts_72;
  assign rport_io_ins_73 = regOuts_73;
  assign rport_io_ins_74 = regOuts_74;
  assign rport_io_ins_75 = regOuts_75;
  assign rport_io_ins_76 = regOuts_76;
  assign rport_io_ins_77 = regOuts_77;
  assign rport_io_ins_78 = regOuts_78;
  assign rport_io_ins_79 = regOuts_79;
  assign rport_io_ins_80 = regOuts_80;
  assign rport_io_ins_81 = regOuts_81;
  assign rport_io_ins_82 = regOuts_82;
  assign rport_io_ins_83 = regOuts_83;
  assign rport_io_ins_84 = regOuts_84;
  assign rport_io_ins_85 = regOuts_85;
  assign rport_io_ins_86 = regOuts_86;
  assign rport_io_ins_87 = regOuts_87;
  assign rport_io_ins_88 = regOuts_88;
  assign rport_io_ins_89 = regOuts_89;
  assign rport_io_ins_90 = regOuts_90;
  assign rport_io_ins_91 = regOuts_91;
  assign rport_io_ins_92 = regOuts_92;
  assign rport_io_ins_93 = regOuts_93;
  assign rport_io_ins_94 = regOuts_94;
  assign rport_io_ins_95 = regOuts_95;
  assign rport_io_ins_96 = regOuts_96;
  assign rport_io_ins_97 = regOuts_97;
  assign rport_io_ins_98 = regOuts_98;
  assign rport_io_ins_99 = regOuts_99;
  assign rport_io_ins_100 = regOuts_100;
  assign rport_io_ins_101 = regOuts_101;
  assign rport_io_ins_102 = regOuts_102;
  assign rport_io_ins_103 = regOuts_103;
  assign rport_io_ins_104 = regOuts_104;
  assign rport_io_ins_105 = regOuts_105;
  assign rport_io_ins_106 = regOuts_106;
  assign rport_io_ins_107 = regOuts_107;
  assign rport_io_ins_108 = regOuts_108;
  assign rport_io_ins_109 = regOuts_109;
  assign rport_io_ins_110 = regOuts_110;
  assign rport_io_ins_111 = regOuts_111;
  assign rport_io_ins_112 = regOuts_112;
  assign rport_io_ins_113 = regOuts_113;
  assign rport_io_ins_114 = regOuts_114;
  assign rport_io_ins_115 = regOuts_115;
  assign rport_io_ins_116 = regOuts_116;
  assign rport_io_ins_117 = regOuts_117;
  assign rport_io_ins_118 = regOuts_118;
  assign rport_io_ins_119 = regOuts_119;
  assign rport_io_ins_120 = regOuts_120;
  assign rport_io_ins_121 = regOuts_121;
  assign rport_io_ins_122 = regOuts_122;
  assign rport_io_ins_123 = regOuts_123;
  assign rport_io_ins_124 = regOuts_124;
  assign rport_io_ins_125 = regOuts_125;
  assign rport_io_ins_126 = regOuts_126;
  assign rport_io_ins_127 = regOuts_127;
  assign rport_io_ins_128 = regOuts_128;
  assign rport_io_ins_129 = regOuts_129;
  assign rport_io_ins_130 = regOuts_130;
  assign rport_io_ins_131 = regOuts_131;
  assign rport_io_ins_132 = regOuts_132;
  assign rport_io_ins_133 = regOuts_133;
  assign rport_io_ins_134 = regOuts_134;
  assign rport_io_ins_135 = regOuts_135;
  assign rport_io_ins_136 = regOuts_136;
  assign rport_io_ins_137 = regOuts_137;
  assign rport_io_ins_138 = regOuts_138;
  assign rport_io_ins_139 = regOuts_139;
  assign rport_io_ins_140 = regOuts_140;
  assign rport_io_ins_141 = regOuts_141;
  assign rport_io_ins_142 = regOuts_142;
  assign rport_io_ins_143 = regOuts_143;
  assign rport_io_ins_144 = regOuts_144;
  assign rport_io_ins_145 = regOuts_145;
  assign rport_io_ins_146 = regOuts_146;
  assign rport_io_ins_147 = regOuts_147;
  assign rport_io_ins_148 = regOuts_148;
  assign rport_io_ins_149 = regOuts_149;
  assign rport_io_ins_150 = regOuts_150;
  assign rport_io_ins_151 = regOuts_151;
  assign rport_io_ins_152 = regOuts_152;
  assign rport_io_ins_153 = regOuts_153;
  assign rport_io_ins_154 = regOuts_154;
  assign rport_io_ins_155 = regOuts_155;
  assign rport_io_ins_156 = regOuts_156;
  assign rport_io_ins_157 = regOuts_157;
  assign rport_io_ins_158 = regOuts_158;
  assign rport_io_ins_159 = regOuts_159;
  assign rport_io_ins_160 = regOuts_160;
  assign rport_io_ins_161 = regOuts_161;
  assign rport_io_ins_162 = regOuts_162;
  assign rport_io_ins_163 = regOuts_163;
  assign rport_io_ins_164 = regOuts_164;
  assign rport_io_ins_165 = regOuts_165;
  assign rport_io_ins_166 = regOuts_166;
  assign rport_io_ins_167 = regOuts_167;
  assign rport_io_ins_168 = regOuts_168;
  assign rport_io_ins_169 = regOuts_169;
  assign rport_io_ins_170 = regOuts_170;
  assign rport_io_ins_171 = regOuts_171;
  assign rport_io_ins_172 = regOuts_172;
  assign rport_io_ins_173 = regOuts_173;
  assign rport_io_ins_174 = regOuts_174;
  assign rport_io_ins_175 = regOuts_175;
  assign rport_io_ins_176 = regOuts_176;
  assign rport_io_ins_177 = regOuts_177;
  assign rport_io_ins_178 = regOuts_178;
  assign rport_io_ins_179 = regOuts_179;
  assign rport_io_ins_180 = regOuts_180;
  assign rport_io_ins_181 = regOuts_181;
  assign rport_io_ins_182 = regOuts_182;
  assign rport_io_ins_183 = regOuts_183;
  assign rport_io_ins_184 = regOuts_184;
  assign rport_io_ins_185 = regOuts_185;
  assign rport_io_ins_186 = regOuts_186;
  assign rport_io_ins_187 = regOuts_187;
  assign rport_io_ins_188 = regOuts_188;
  assign rport_io_ins_189 = regOuts_189;
  assign rport_io_ins_190 = regOuts_190;
  assign rport_io_ins_191 = regOuts_191;
  assign rport_io_ins_192 = regOuts_192;
  assign rport_io_ins_193 = regOuts_193;
  assign rport_io_ins_194 = regOuts_194;
  assign rport_io_ins_195 = regOuts_195;
  assign rport_io_ins_196 = regOuts_196;
  assign rport_io_ins_197 = regOuts_197;
  assign rport_io_ins_198 = regOuts_198;
  assign rport_io_ins_199 = regOuts_199;
  assign rport_io_ins_200 = regOuts_200;
  assign rport_io_ins_201 = regOuts_201;
  assign rport_io_ins_202 = regOuts_202;
  assign rport_io_ins_203 = regOuts_203;
  assign rport_io_ins_204 = regOuts_204;
  assign rport_io_ins_205 = regOuts_205;
  assign rport_io_ins_206 = regOuts_206;
  assign rport_io_ins_207 = regOuts_207;
  assign rport_io_ins_208 = regOuts_208;
  assign rport_io_ins_209 = regOuts_209;
  assign rport_io_ins_210 = regOuts_210;
  assign rport_io_ins_211 = regOuts_211;
  assign rport_io_ins_212 = regOuts_212;
  assign rport_io_ins_213 = regOuts_213;
  assign rport_io_ins_214 = regOuts_214;
  assign rport_io_ins_215 = regOuts_215;
  assign rport_io_ins_216 = regOuts_216;
  assign rport_io_ins_217 = regOuts_217;
  assign rport_io_ins_218 = regOuts_218;
  assign rport_io_ins_219 = regOuts_219;
  assign rport_io_ins_220 = regOuts_220;
  assign rport_io_ins_221 = regOuts_221;
  assign rport_io_ins_222 = regOuts_222;
  assign rport_io_ins_223 = regOuts_223;
  assign rport_io_ins_224 = regOuts_224;
  assign rport_io_ins_225 = regOuts_225;
  assign rport_io_ins_226 = regOuts_226;
  assign rport_io_ins_227 = regOuts_227;
  assign rport_io_ins_228 = regOuts_228;
  assign rport_io_ins_229 = regOuts_229;
  assign rport_io_ins_230 = regOuts_230;
  assign rport_io_ins_231 = regOuts_231;
  assign rport_io_ins_232 = regOuts_232;
  assign rport_io_ins_233 = regOuts_233;
  assign rport_io_ins_234 = regOuts_234;
  assign rport_io_ins_235 = regOuts_235;
  assign rport_io_sel = io_raddr;
  assign regOuts_0 = regs_0_io_out;
  assign regOuts_1 = regs_1_io_out;
  assign regOuts_2 = regs_2_io_out;
  assign regOuts_3 = regs_3_io_out;
  assign regOuts_4 = regs_4_io_out;
  assign regOuts_5 = regs_5_io_out;
  assign regOuts_6 = regs_6_io_out;
  assign regOuts_7 = regs_7_io_out;
  assign regOuts_8 = regs_8_io_out;
  assign regOuts_9 = regs_9_io_out;
  assign regOuts_10 = regs_10_io_out;
  assign regOuts_11 = regs_11_io_out;
  assign regOuts_12 = regs_12_io_out;
  assign regOuts_13 = regs_13_io_out;
  assign regOuts_14 = regs_14_io_out;
  assign regOuts_15 = regs_15_io_out;
  assign regOuts_16 = regs_16_io_out;
  assign regOuts_17 = regs_17_io_out;
  assign regOuts_18 = regs_18_io_out;
  assign regOuts_19 = regs_19_io_out;
  assign regOuts_20 = regs_20_io_out;
  assign regOuts_21 = regs_21_io_out;
  assign regOuts_22 = regs_22_io_out;
  assign regOuts_23 = regs_23_io_out;
  assign regOuts_24 = regs_24_io_out;
  assign regOuts_25 = regs_25_io_out;
  assign regOuts_26 = regs_26_io_out;
  assign regOuts_27 = regs_27_io_out;
  assign regOuts_28 = regs_28_io_out;
  assign regOuts_29 = regs_29_io_out;
  assign regOuts_30 = regs_30_io_out;
  assign regOuts_31 = regs_31_io_out;
  assign regOuts_32 = regs_32_io_out;
  assign regOuts_33 = regs_33_io_out;
  assign regOuts_34 = regs_34_io_out;
  assign regOuts_35 = regs_35_io_out;
  assign regOuts_36 = regs_36_io_out;
  assign regOuts_37 = regs_37_io_out;
  assign regOuts_38 = regs_38_io_out;
  assign regOuts_39 = regs_39_io_out;
  assign regOuts_40 = regs_40_io_out;
  assign regOuts_41 = regs_41_io_out;
  assign regOuts_42 = regs_42_io_out;
  assign regOuts_43 = regs_43_io_out;
  assign regOuts_44 = regs_44_io_out;
  assign regOuts_45 = regs_45_io_out;
  assign regOuts_46 = regs_46_io_out;
  assign regOuts_47 = regs_47_io_out;
  assign regOuts_48 = regs_48_io_out;
  assign regOuts_49 = regs_49_io_out;
  assign regOuts_50 = regs_50_io_out;
  assign regOuts_51 = regs_51_io_out;
  assign regOuts_52 = regs_52_io_out;
  assign regOuts_53 = regs_53_io_out;
  assign regOuts_54 = regs_54_io_out;
  assign regOuts_55 = regs_55_io_out;
  assign regOuts_56 = regs_56_io_out;
  assign regOuts_57 = regs_57_io_out;
  assign regOuts_58 = regs_58_io_out;
  assign regOuts_59 = regs_59_io_out;
  assign regOuts_60 = regs_60_io_out;
  assign regOuts_61 = regs_61_io_out;
  assign regOuts_62 = regs_62_io_out;
  assign regOuts_63 = regs_63_io_out;
  assign regOuts_64 = regs_64_io_out;
  assign regOuts_65 = regs_65_io_out;
  assign regOuts_66 = regs_66_io_out;
  assign regOuts_67 = regs_67_io_out;
  assign regOuts_68 = regs_68_io_out;
  assign regOuts_69 = regs_69_io_out;
  assign regOuts_70 = regs_70_io_out;
  assign regOuts_71 = regs_71_io_out;
  assign regOuts_72 = regs_72_io_out;
  assign regOuts_73 = regs_73_io_out;
  assign regOuts_74 = regs_74_io_out;
  assign regOuts_75 = regs_75_io_out;
  assign regOuts_76 = regs_76_io_out;
  assign regOuts_77 = regs_77_io_out;
  assign regOuts_78 = regs_78_io_out;
  assign regOuts_79 = regs_79_io_out;
  assign regOuts_80 = regs_80_io_out;
  assign regOuts_81 = regs_81_io_out;
  assign regOuts_82 = regs_82_io_out;
  assign regOuts_83 = regs_83_io_out;
  assign regOuts_84 = regs_84_io_out;
  assign regOuts_85 = regs_85_io_out;
  assign regOuts_86 = regs_86_io_out;
  assign regOuts_87 = regs_87_io_out;
  assign regOuts_88 = regs_88_io_out;
  assign regOuts_89 = regs_89_io_out;
  assign regOuts_90 = regs_90_io_out;
  assign regOuts_91 = regs_91_io_out;
  assign regOuts_92 = regs_92_io_out;
  assign regOuts_93 = regs_93_io_out;
  assign regOuts_94 = regs_94_io_out;
  assign regOuts_95 = regs_95_io_out;
  assign regOuts_96 = regs_96_io_out;
  assign regOuts_97 = regs_97_io_out;
  assign regOuts_98 = regs_98_io_out;
  assign regOuts_99 = regs_99_io_out;
  assign regOuts_100 = regs_100_io_out;
  assign regOuts_101 = regs_101_io_out;
  assign regOuts_102 = regs_102_io_out;
  assign regOuts_103 = regs_103_io_out;
  assign regOuts_104 = regs_104_io_out;
  assign regOuts_105 = regs_105_io_out;
  assign regOuts_106 = regs_106_io_out;
  assign regOuts_107 = regs_107_io_out;
  assign regOuts_108 = regs_108_io_out;
  assign regOuts_109 = regs_109_io_out;
  assign regOuts_110 = regs_110_io_out;
  assign regOuts_111 = regs_111_io_out;
  assign regOuts_112 = regs_112_io_out;
  assign regOuts_113 = regs_113_io_out;
  assign regOuts_114 = regs_114_io_out;
  assign regOuts_115 = regs_115_io_out;
  assign regOuts_116 = regs_116_io_out;
  assign regOuts_117 = regs_117_io_out;
  assign regOuts_118 = regs_118_io_out;
  assign regOuts_119 = regs_119_io_out;
  assign regOuts_120 = regs_120_io_out;
  assign regOuts_121 = regs_121_io_out;
  assign regOuts_122 = regs_122_io_out;
  assign regOuts_123 = regs_123_io_out;
  assign regOuts_124 = regs_124_io_out;
  assign regOuts_125 = regs_125_io_out;
  assign regOuts_126 = regs_126_io_out;
  assign regOuts_127 = regs_127_io_out;
  assign regOuts_128 = regs_128_io_out;
  assign regOuts_129 = regs_129_io_out;
  assign regOuts_130 = regs_130_io_out;
  assign regOuts_131 = regs_131_io_out;
  assign regOuts_132 = regs_132_io_out;
  assign regOuts_133 = regs_133_io_out;
  assign regOuts_134 = regs_134_io_out;
  assign regOuts_135 = regs_135_io_out;
  assign regOuts_136 = regs_136_io_out;
  assign regOuts_137 = regs_137_io_out;
  assign regOuts_138 = regs_138_io_out;
  assign regOuts_139 = regs_139_io_out;
  assign regOuts_140 = regs_140_io_out;
  assign regOuts_141 = regs_141_io_out;
  assign regOuts_142 = regs_142_io_out;
  assign regOuts_143 = regs_143_io_out;
  assign regOuts_144 = regs_144_io_out;
  assign regOuts_145 = regs_145_io_out;
  assign regOuts_146 = regs_146_io_out;
  assign regOuts_147 = regs_147_io_out;
  assign regOuts_148 = regs_148_io_out;
  assign regOuts_149 = regs_149_io_out;
  assign regOuts_150 = regs_150_io_out;
  assign regOuts_151 = regs_151_io_out;
  assign regOuts_152 = regs_152_io_out;
  assign regOuts_153 = regs_153_io_out;
  assign regOuts_154 = regs_154_io_out;
  assign regOuts_155 = regs_155_io_out;
  assign regOuts_156 = regs_156_io_out;
  assign regOuts_157 = regs_157_io_out;
  assign regOuts_158 = regs_158_io_out;
  assign regOuts_159 = regs_159_io_out;
  assign regOuts_160 = regs_160_io_out;
  assign regOuts_161 = regs_161_io_out;
  assign regOuts_162 = regs_162_io_out;
  assign regOuts_163 = regs_163_io_out;
  assign regOuts_164 = regs_164_io_out;
  assign regOuts_165 = regs_165_io_out;
  assign regOuts_166 = regs_166_io_out;
  assign regOuts_167 = regs_167_io_out;
  assign regOuts_168 = regs_168_io_out;
  assign regOuts_169 = regs_169_io_out;
  assign regOuts_170 = regs_170_io_out;
  assign regOuts_171 = regs_171_io_out;
  assign regOuts_172 = regs_172_io_out;
  assign regOuts_173 = regs_173_io_out;
  assign regOuts_174 = regs_174_io_out;
  assign regOuts_175 = regs_175_io_out;
  assign regOuts_176 = regs_176_io_out;
  assign regOuts_177 = regs_177_io_out;
  assign regOuts_178 = regs_178_io_out;
  assign regOuts_179 = regs_179_io_out;
  assign regOuts_180 = regs_180_io_out;
  assign regOuts_181 = regs_181_io_out;
  assign regOuts_182 = regs_182_io_out;
  assign regOuts_183 = regs_183_io_out;
  assign regOuts_184 = regs_184_io_out;
  assign regOuts_185 = regs_185_io_out;
  assign regOuts_186 = regs_186_io_out;
  assign regOuts_187 = regs_187_io_out;
  assign regOuts_188 = regs_188_io_out;
  assign regOuts_189 = regs_189_io_out;
  assign regOuts_190 = regs_190_io_out;
  assign regOuts_191 = regs_191_io_out;
  assign regOuts_192 = regs_192_io_out;
  assign regOuts_193 = regs_193_io_out;
  assign regOuts_194 = regs_194_io_out;
  assign regOuts_195 = regs_195_io_out;
  assign regOuts_196 = regs_196_io_out;
  assign regOuts_197 = regs_197_io_out;
  assign regOuts_198 = regs_198_io_out;
  assign regOuts_199 = regs_199_io_out;
  assign regOuts_200 = regs_200_io_out;
  assign regOuts_201 = regs_201_io_out;
  assign regOuts_202 = regs_202_io_out;
  assign regOuts_203 = regs_203_io_out;
  assign regOuts_204 = regs_204_io_out;
  assign regOuts_205 = regs_205_io_out;
  assign regOuts_206 = regs_206_io_out;
  assign regOuts_207 = regs_207_io_out;
  assign regOuts_208 = regs_208_io_out;
  assign regOuts_209 = regs_209_io_out;
  assign regOuts_210 = regs_210_io_out;
  assign regOuts_211 = regs_211_io_out;
  assign regOuts_212 = regs_212_io_out;
  assign regOuts_213 = regs_213_io_out;
  assign regOuts_214 = regs_214_io_out;
  assign regOuts_215 = regs_215_io_out;
  assign regOuts_216 = regs_216_io_out;
  assign regOuts_217 = regs_217_io_out;
  assign regOuts_218 = regs_218_io_out;
  assign regOuts_219 = regs_219_io_out;
  assign regOuts_220 = regs_220_io_out;
  assign regOuts_221 = regs_221_io_out;
  assign regOuts_222 = regs_222_io_out;
  assign regOuts_223 = regs_223_io_out;
  assign regOuts_224 = regs_224_io_out;
  assign regOuts_225 = regs_225_io_out;
  assign regOuts_226 = regs_226_io_out;
  assign regOuts_227 = regs_227_io_out;
  assign regOuts_228 = regs_228_io_out;
  assign regOuts_229 = regs_229_io_out;
  assign regOuts_230 = regs_230_io_out;
  assign regOuts_231 = regs_231_io_out;
  assign regOuts_232 = regs_232_io_out;
  assign regOuts_233 = regs_233_io_out;
  assign regOuts_234 = regs_234_io_out;
  assign regOuts_235 = regs_235_io_out;
  assign _T_2390_0 = regOuts_0;
  assign _T_2390_1 = regOuts_1;
  assign _T_2390_2 = regOuts_2;
endmodule
module Fringe(
  input         clock,
  input         reset,
  input  [31:0] io_raddr,
  input         io_wen,
  input  [31:0] io_waddr,
  input  [63:0] io_wdata,
  output [63:0] io_rdata,
  output        io_enable,
  input         io_done,
  output [63:0] io_argIns_0,
  input         io_argOuts_0_valid,
  input  [63:0] io_argOuts_0_bits
);
  wire  mags_0_clock;
  wire  mags_0_reset;
  wire  mags_0_io_enable;
  wire [31:0] mags_0_io_debugSignals_0;
  wire [31:0] mags_0_io_debugSignals_1;
  wire [31:0] mags_0_io_debugSignals_2;
  wire [31:0] mags_0_io_debugSignals_3;
  wire [31:0] mags_0_io_debugSignals_4;
  wire [31:0] mags_0_io_debugSignals_5;
  wire [31:0] mags_0_io_debugSignals_6;
  wire [31:0] mags_0_io_debugSignals_7;
  wire [31:0] mags_0_io_debugSignals_8;
  wire [31:0] mags_0_io_debugSignals_9;
  wire [31:0] mags_0_io_debugSignals_10;
  wire [31:0] mags_0_io_debugSignals_11;
  wire [31:0] mags_0_io_debugSignals_12;
  wire [31:0] mags_0_io_debugSignals_13;
  wire [31:0] mags_0_io_debugSignals_14;
  wire [31:0] mags_0_io_debugSignals_15;
  wire [31:0] mags_0_io_debugSignals_16;
  wire [31:0] mags_0_io_debugSignals_17;
  wire [31:0] mags_0_io_debugSignals_18;
  wire [31:0] mags_0_io_debugSignals_19;
  wire [31:0] mags_0_io_debugSignals_20;
  wire [31:0] mags_0_io_debugSignals_21;
  wire [31:0] mags_0_io_debugSignals_22;
  wire [31:0] mags_0_io_debugSignals_23;
  wire [31:0] mags_0_io_debugSignals_24;
  wire [31:0] mags_0_io_debugSignals_25;
  wire [31:0] mags_0_io_debugSignals_26;
  wire [31:0] mags_0_io_debugSignals_27;
  wire [31:0] mags_0_io_debugSignals_28;
  wire [31:0] mags_0_io_debugSignals_29;
  wire [31:0] mags_0_io_debugSignals_30;
  wire [31:0] mags_0_io_debugSignals_31;
  wire [31:0] mags_0_io_debugSignals_32;
  wire [31:0] mags_0_io_debugSignals_33;
  wire [31:0] mags_0_io_debugSignals_34;
  wire [31:0] mags_0_io_debugSignals_35;
  wire [31:0] mags_0_io_debugSignals_36;
  wire [31:0] mags_0_io_debugSignals_37;
  wire [31:0] mags_0_io_debugSignals_38;
  wire [31:0] mags_0_io_debugSignals_39;
  wire [31:0] mags_0_io_debugSignals_40;
  wire [31:0] mags_0_io_debugSignals_41;
  wire [31:0] mags_0_io_debugSignals_42;
  wire [31:0] mags_0_io_debugSignals_43;
  wire [31:0] mags_0_io_debugSignals_44;
  wire [31:0] mags_0_io_debugSignals_45;
  wire [31:0] mags_0_io_debugSignals_46;
  wire [31:0] mags_0_io_debugSignals_47;
  wire [31:0] mags_0_io_debugSignals_48;
  wire [31:0] mags_0_io_debugSignals_49;
  wire [31:0] mags_0_io_debugSignals_50;
  wire [31:0] mags_0_io_debugSignals_51;
  wire [31:0] mags_0_io_debugSignals_52;
  wire [31:0] mags_0_io_debugSignals_53;
  wire [31:0] mags_0_io_debugSignals_54;
  wire [31:0] mags_0_io_debugSignals_55;
  wire [31:0] mags_0_io_debugSignals_56;
  wire [31:0] mags_0_io_debugSignals_57;
  wire [31:0] mags_0_io_debugSignals_58;
  wire  mags_0_io_dram_rresp_ready;
  wire  regs_clock;
  wire  regs_reset;
  wire [7:0] regs_io_raddr;
  wire  regs_io_wen;
  wire [7:0] regs_io_waddr;
  wire [63:0] regs_io_wdata;
  wire [63:0] regs_io_rdata;
  wire [63:0] regs_io_argIns_0;
  wire [63:0] regs_io_argIns_1;
  wire [63:0] regs_io_argIns_2;
  wire  regs_io_argOuts_0_valid;
  wire [63:0] regs_io_argOuts_0_bits;
  wire  regs_io_argOuts_1_valid;
  wire [63:0] regs_io_argOuts_1_bits;
  wire [63:0] regs_io_argOuts_2_bits;
  wire [63:0] regs_io_argOuts_3_bits;
  wire [63:0] regs_io_argOuts_4_bits;
  wire [63:0] regs_io_argOuts_5_bits;
  wire [63:0] regs_io_argOuts_6_bits;
  wire [63:0] regs_io_argOuts_7_bits;
  wire [63:0] regs_io_argOuts_8_bits;
  wire [63:0] regs_io_argOuts_9_bits;
  wire [63:0] regs_io_argOuts_10_bits;
  wire [63:0] regs_io_argOuts_11_bits;
  wire [63:0] regs_io_argOuts_12_bits;
  wire [63:0] regs_io_argOuts_13_bits;
  wire [63:0] regs_io_argOuts_14_bits;
  wire [63:0] regs_io_argOuts_15_bits;
  wire [63:0] regs_io_argOuts_16_bits;
  wire [63:0] regs_io_argOuts_17_bits;
  wire [63:0] regs_io_argOuts_18_bits;
  wire [63:0] regs_io_argOuts_19_bits;
  wire [63:0] regs_io_argOuts_20_bits;
  wire [63:0] regs_io_argOuts_21_bits;
  wire [63:0] regs_io_argOuts_22_bits;
  wire [63:0] regs_io_argOuts_23_bits;
  wire [63:0] regs_io_argOuts_24_bits;
  wire [63:0] regs_io_argOuts_25_bits;
  wire [63:0] regs_io_argOuts_26_bits;
  wire [63:0] regs_io_argOuts_27_bits;
  wire [63:0] regs_io_argOuts_28_bits;
  wire [63:0] regs_io_argOuts_29_bits;
  wire [63:0] regs_io_argOuts_30_bits;
  wire [63:0] regs_io_argOuts_31_bits;
  wire [63:0] regs_io_argOuts_32_bits;
  wire [63:0] regs_io_argOuts_33_bits;
  wire [63:0] regs_io_argOuts_34_bits;
  wire [63:0] regs_io_argOuts_35_bits;
  wire [63:0] regs_io_argOuts_36_bits;
  wire [63:0] regs_io_argOuts_37_bits;
  wire [63:0] regs_io_argOuts_38_bits;
  wire [63:0] regs_io_argOuts_39_bits;
  wire [63:0] regs_io_argOuts_40_bits;
  wire [63:0] regs_io_argOuts_41_bits;
  wire [63:0] regs_io_argOuts_42_bits;
  wire [63:0] regs_io_argOuts_43_bits;
  wire [63:0] regs_io_argOuts_44_bits;
  wire [63:0] regs_io_argOuts_45_bits;
  wire [63:0] regs_io_argOuts_46_bits;
  wire [63:0] regs_io_argOuts_47_bits;
  wire [63:0] regs_io_argOuts_48_bits;
  wire [63:0] regs_io_argOuts_49_bits;
  wire [63:0] regs_io_argOuts_50_bits;
  wire [63:0] regs_io_argOuts_51_bits;
  wire [63:0] regs_io_argOuts_52_bits;
  wire [63:0] regs_io_argOuts_53_bits;
  wire [63:0] regs_io_argOuts_54_bits;
  wire [63:0] regs_io_argOuts_55_bits;
  wire [63:0] regs_io_argOuts_56_bits;
  wire [63:0] regs_io_argOuts_57_bits;
  wire [63:0] regs_io_argOuts_58_bits;
  wire [63:0] regs_io_argOuts_59_bits;
  wire [63:0] regs_io_argOuts_60_bits;
  wire  _T_351;
  wire  _T_352;
  wire  _T_353;
  wire  localEnable;
  wire  timeoutCtr_clock;
  wire  timeoutCtr_reset;
  wire [39:0] timeoutCtr_io_max;
  wire [39:0] timeoutCtr_io_out;
  wire  timeoutCtr_io_enable;
  wire  timeoutCtr_io_saturate;
  wire  timeoutCtr_io_done;
  wire  depulser_clock;
  wire  depulser_reset;
  wire  depulser_io_in;
  wire  depulser_io_rst;
  wire  depulser_io_out;
  wire  _T_358;
  wire [63:0] _T_359;
  wire  status_valid;
  wire [63:0] status_bits;
  wire  _T_369;
  wire  _T_371;
  wire [1:0] _T_372;
  MAGCore mags_0 (
    .clock(mags_0_clock),
    .reset(mags_0_reset),
    .io_enable(mags_0_io_enable),
    .io_debugSignals_0(mags_0_io_debugSignals_0),
    .io_debugSignals_1(mags_0_io_debugSignals_1),
    .io_debugSignals_2(mags_0_io_debugSignals_2),
    .io_debugSignals_3(mags_0_io_debugSignals_3),
    .io_debugSignals_4(mags_0_io_debugSignals_4),
    .io_debugSignals_5(mags_0_io_debugSignals_5),
    .io_debugSignals_6(mags_0_io_debugSignals_6),
    .io_debugSignals_7(mags_0_io_debugSignals_7),
    .io_debugSignals_8(mags_0_io_debugSignals_8),
    .io_debugSignals_9(mags_0_io_debugSignals_9),
    .io_debugSignals_10(mags_0_io_debugSignals_10),
    .io_debugSignals_11(mags_0_io_debugSignals_11),
    .io_debugSignals_12(mags_0_io_debugSignals_12),
    .io_debugSignals_13(mags_0_io_debugSignals_13),
    .io_debugSignals_14(mags_0_io_debugSignals_14),
    .io_debugSignals_15(mags_0_io_debugSignals_15),
    .io_debugSignals_16(mags_0_io_debugSignals_16),
    .io_debugSignals_17(mags_0_io_debugSignals_17),
    .io_debugSignals_18(mags_0_io_debugSignals_18),
    .io_debugSignals_19(mags_0_io_debugSignals_19),
    .io_debugSignals_20(mags_0_io_debugSignals_20),
    .io_debugSignals_21(mags_0_io_debugSignals_21),
    .io_debugSignals_22(mags_0_io_debugSignals_22),
    .io_debugSignals_23(mags_0_io_debugSignals_23),
    .io_debugSignals_24(mags_0_io_debugSignals_24),
    .io_debugSignals_25(mags_0_io_debugSignals_25),
    .io_debugSignals_26(mags_0_io_debugSignals_26),
    .io_debugSignals_27(mags_0_io_debugSignals_27),
    .io_debugSignals_28(mags_0_io_debugSignals_28),
    .io_debugSignals_29(mags_0_io_debugSignals_29),
    .io_debugSignals_30(mags_0_io_debugSignals_30),
    .io_debugSignals_31(mags_0_io_debugSignals_31),
    .io_debugSignals_32(mags_0_io_debugSignals_32),
    .io_debugSignals_33(mags_0_io_debugSignals_33),
    .io_debugSignals_34(mags_0_io_debugSignals_34),
    .io_debugSignals_35(mags_0_io_debugSignals_35),
    .io_debugSignals_36(mags_0_io_debugSignals_36),
    .io_debugSignals_37(mags_0_io_debugSignals_37),
    .io_debugSignals_38(mags_0_io_debugSignals_38),
    .io_debugSignals_39(mags_0_io_debugSignals_39),
    .io_debugSignals_40(mags_0_io_debugSignals_40),
    .io_debugSignals_41(mags_0_io_debugSignals_41),
    .io_debugSignals_42(mags_0_io_debugSignals_42),
    .io_debugSignals_43(mags_0_io_debugSignals_43),
    .io_debugSignals_44(mags_0_io_debugSignals_44),
    .io_debugSignals_45(mags_0_io_debugSignals_45),
    .io_debugSignals_46(mags_0_io_debugSignals_46),
    .io_debugSignals_47(mags_0_io_debugSignals_47),
    .io_debugSignals_48(mags_0_io_debugSignals_48),
    .io_debugSignals_49(mags_0_io_debugSignals_49),
    .io_debugSignals_50(mags_0_io_debugSignals_50),
    .io_debugSignals_51(mags_0_io_debugSignals_51),
    .io_debugSignals_52(mags_0_io_debugSignals_52),
    .io_debugSignals_53(mags_0_io_debugSignals_53),
    .io_debugSignals_54(mags_0_io_debugSignals_54),
    .io_debugSignals_55(mags_0_io_debugSignals_55),
    .io_debugSignals_56(mags_0_io_debugSignals_56),
    .io_debugSignals_57(mags_0_io_debugSignals_57),
    .io_debugSignals_58(mags_0_io_debugSignals_58),
    .io_dram_rresp_ready(mags_0_io_dram_rresp_ready)
  );
  RegFile regs (
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits),
    .io_argOuts_2_bits(regs_io_argOuts_2_bits),
    .io_argOuts_3_bits(regs_io_argOuts_3_bits),
    .io_argOuts_4_bits(regs_io_argOuts_4_bits),
    .io_argOuts_5_bits(regs_io_argOuts_5_bits),
    .io_argOuts_6_bits(regs_io_argOuts_6_bits),
    .io_argOuts_7_bits(regs_io_argOuts_7_bits),
    .io_argOuts_8_bits(regs_io_argOuts_8_bits),
    .io_argOuts_9_bits(regs_io_argOuts_9_bits),
    .io_argOuts_10_bits(regs_io_argOuts_10_bits),
    .io_argOuts_11_bits(regs_io_argOuts_11_bits),
    .io_argOuts_12_bits(regs_io_argOuts_12_bits),
    .io_argOuts_13_bits(regs_io_argOuts_13_bits),
    .io_argOuts_14_bits(regs_io_argOuts_14_bits),
    .io_argOuts_15_bits(regs_io_argOuts_15_bits),
    .io_argOuts_16_bits(regs_io_argOuts_16_bits),
    .io_argOuts_17_bits(regs_io_argOuts_17_bits),
    .io_argOuts_18_bits(regs_io_argOuts_18_bits),
    .io_argOuts_19_bits(regs_io_argOuts_19_bits),
    .io_argOuts_20_bits(regs_io_argOuts_20_bits),
    .io_argOuts_21_bits(regs_io_argOuts_21_bits),
    .io_argOuts_22_bits(regs_io_argOuts_22_bits),
    .io_argOuts_23_bits(regs_io_argOuts_23_bits),
    .io_argOuts_24_bits(regs_io_argOuts_24_bits),
    .io_argOuts_25_bits(regs_io_argOuts_25_bits),
    .io_argOuts_26_bits(regs_io_argOuts_26_bits),
    .io_argOuts_27_bits(regs_io_argOuts_27_bits),
    .io_argOuts_28_bits(regs_io_argOuts_28_bits),
    .io_argOuts_29_bits(regs_io_argOuts_29_bits),
    .io_argOuts_30_bits(regs_io_argOuts_30_bits),
    .io_argOuts_31_bits(regs_io_argOuts_31_bits),
    .io_argOuts_32_bits(regs_io_argOuts_32_bits),
    .io_argOuts_33_bits(regs_io_argOuts_33_bits),
    .io_argOuts_34_bits(regs_io_argOuts_34_bits),
    .io_argOuts_35_bits(regs_io_argOuts_35_bits),
    .io_argOuts_36_bits(regs_io_argOuts_36_bits),
    .io_argOuts_37_bits(regs_io_argOuts_37_bits),
    .io_argOuts_38_bits(regs_io_argOuts_38_bits),
    .io_argOuts_39_bits(regs_io_argOuts_39_bits),
    .io_argOuts_40_bits(regs_io_argOuts_40_bits),
    .io_argOuts_41_bits(regs_io_argOuts_41_bits),
    .io_argOuts_42_bits(regs_io_argOuts_42_bits),
    .io_argOuts_43_bits(regs_io_argOuts_43_bits),
    .io_argOuts_44_bits(regs_io_argOuts_44_bits),
    .io_argOuts_45_bits(regs_io_argOuts_45_bits),
    .io_argOuts_46_bits(regs_io_argOuts_46_bits),
    .io_argOuts_47_bits(regs_io_argOuts_47_bits),
    .io_argOuts_48_bits(regs_io_argOuts_48_bits),
    .io_argOuts_49_bits(regs_io_argOuts_49_bits),
    .io_argOuts_50_bits(regs_io_argOuts_50_bits),
    .io_argOuts_51_bits(regs_io_argOuts_51_bits),
    .io_argOuts_52_bits(regs_io_argOuts_52_bits),
    .io_argOuts_53_bits(regs_io_argOuts_53_bits),
    .io_argOuts_54_bits(regs_io_argOuts_54_bits),
    .io_argOuts_55_bits(regs_io_argOuts_55_bits),
    .io_argOuts_56_bits(regs_io_argOuts_56_bits),
    .io_argOuts_57_bits(regs_io_argOuts_57_bits),
    .io_argOuts_58_bits(regs_io_argOuts_58_bits),
    .io_argOuts_59_bits(regs_io_argOuts_59_bits),
    .io_argOuts_60_bits(regs_io_argOuts_60_bits)
  );
  Counter_19 timeoutCtr (
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_max(timeoutCtr_io_max),
    .io_out(timeoutCtr_io_out),
    .io_enable(timeoutCtr_io_enable),
    .io_saturate(timeoutCtr_io_saturate),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser (
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_351 = regs_io_argIns_0[0];
  assign _T_352 = regs_io_argIns_1[0];
  assign _T_353 = ~ _T_352;
  assign localEnable = _T_351 & _T_353;
  assign _T_358 = io_done | timeoutCtr_io_done;
  assign _T_359 = ~ regs_io_argIns_0;
  assign _T_369 = _T_351 & timeoutCtr_io_done;
  assign _T_371 = _T_351 & depulser_io_out;
  assign _T_372 = {_T_369,_T_371};
  assign io_rdata = regs_io_rdata;
  assign io_enable = localEnable;
  assign io_argIns_0 = regs_io_argIns_2;
  assign mags_0_io_enable = localEnable;
  assign mags_0_clock = clock;
  assign mags_0_reset = reset;
  assign regs_io_raddr = io_raddr[7:0];
  assign regs_io_wen = io_wen;
  assign regs_io_waddr = io_waddr[7:0];
  assign regs_io_wdata = io_wdata;
  assign regs_io_argOuts_0_valid = status_valid;
  assign regs_io_argOuts_0_bits = status_bits;
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid;
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits;
  assign regs_io_argOuts_2_bits = {{32'd0}, mags_0_io_debugSignals_0};
  assign regs_io_argOuts_3_bits = {{32'd0}, mags_0_io_debugSignals_1};
  assign regs_io_argOuts_4_bits = {{32'd0}, mags_0_io_debugSignals_2};
  assign regs_io_argOuts_5_bits = {{32'd0}, mags_0_io_debugSignals_3};
  assign regs_io_argOuts_6_bits = {{32'd0}, mags_0_io_debugSignals_4};
  assign regs_io_argOuts_7_bits = {{32'd0}, mags_0_io_debugSignals_5};
  assign regs_io_argOuts_8_bits = {{32'd0}, mags_0_io_debugSignals_6};
  assign regs_io_argOuts_9_bits = {{32'd0}, mags_0_io_debugSignals_7};
  assign regs_io_argOuts_10_bits = {{32'd0}, mags_0_io_debugSignals_8};
  assign regs_io_argOuts_11_bits = {{32'd0}, mags_0_io_debugSignals_9};
  assign regs_io_argOuts_12_bits = {{32'd0}, mags_0_io_debugSignals_10};
  assign regs_io_argOuts_13_bits = {{32'd0}, mags_0_io_debugSignals_11};
  assign regs_io_argOuts_14_bits = {{32'd0}, mags_0_io_debugSignals_12};
  assign regs_io_argOuts_15_bits = {{32'd0}, mags_0_io_debugSignals_13};
  assign regs_io_argOuts_16_bits = {{32'd0}, mags_0_io_debugSignals_14};
  assign regs_io_argOuts_17_bits = {{32'd0}, mags_0_io_debugSignals_15};
  assign regs_io_argOuts_18_bits = {{32'd0}, mags_0_io_debugSignals_16};
  assign regs_io_argOuts_19_bits = {{32'd0}, mags_0_io_debugSignals_17};
  assign regs_io_argOuts_20_bits = {{32'd0}, mags_0_io_debugSignals_18};
  assign regs_io_argOuts_21_bits = {{32'd0}, mags_0_io_debugSignals_19};
  assign regs_io_argOuts_22_bits = {{32'd0}, mags_0_io_debugSignals_20};
  assign regs_io_argOuts_23_bits = {{32'd0}, mags_0_io_debugSignals_21};
  assign regs_io_argOuts_24_bits = {{32'd0}, mags_0_io_debugSignals_22};
  assign regs_io_argOuts_25_bits = {{32'd0}, mags_0_io_debugSignals_23};
  assign regs_io_argOuts_26_bits = {{32'd0}, mags_0_io_debugSignals_24};
  assign regs_io_argOuts_27_bits = {{32'd0}, mags_0_io_debugSignals_25};
  assign regs_io_argOuts_28_bits = {{32'd0}, mags_0_io_debugSignals_26};
  assign regs_io_argOuts_29_bits = {{32'd0}, mags_0_io_debugSignals_27};
  assign regs_io_argOuts_30_bits = {{32'd0}, mags_0_io_debugSignals_28};
  assign regs_io_argOuts_31_bits = {{32'd0}, mags_0_io_debugSignals_29};
  assign regs_io_argOuts_32_bits = {{32'd0}, mags_0_io_debugSignals_30};
  assign regs_io_argOuts_33_bits = {{32'd0}, mags_0_io_debugSignals_31};
  assign regs_io_argOuts_34_bits = {{32'd0}, mags_0_io_debugSignals_32};
  assign regs_io_argOuts_35_bits = {{32'd0}, mags_0_io_debugSignals_33};
  assign regs_io_argOuts_36_bits = {{32'd0}, mags_0_io_debugSignals_34};
  assign regs_io_argOuts_37_bits = {{32'd0}, mags_0_io_debugSignals_35};
  assign regs_io_argOuts_38_bits = {{32'd0}, mags_0_io_debugSignals_36};
  assign regs_io_argOuts_39_bits = {{32'd0}, mags_0_io_debugSignals_37};
  assign regs_io_argOuts_40_bits = {{32'd0}, mags_0_io_debugSignals_38};
  assign regs_io_argOuts_41_bits = {{32'd0}, mags_0_io_debugSignals_39};
  assign regs_io_argOuts_42_bits = {{32'd0}, mags_0_io_debugSignals_40};
  assign regs_io_argOuts_43_bits = {{32'd0}, mags_0_io_debugSignals_41};
  assign regs_io_argOuts_44_bits = {{32'd0}, mags_0_io_debugSignals_42};
  assign regs_io_argOuts_45_bits = {{32'd0}, mags_0_io_debugSignals_43};
  assign regs_io_argOuts_46_bits = {{32'd0}, mags_0_io_debugSignals_44};
  assign regs_io_argOuts_47_bits = {{32'd0}, mags_0_io_debugSignals_45};
  assign regs_io_argOuts_48_bits = {{32'd0}, mags_0_io_debugSignals_46};
  assign regs_io_argOuts_49_bits = {{32'd0}, mags_0_io_debugSignals_47};
  assign regs_io_argOuts_50_bits = {{32'd0}, mags_0_io_debugSignals_48};
  assign regs_io_argOuts_51_bits = {{32'd0}, mags_0_io_debugSignals_49};
  assign regs_io_argOuts_52_bits = {{32'd0}, mags_0_io_debugSignals_50};
  assign regs_io_argOuts_53_bits = {{32'd0}, mags_0_io_debugSignals_51};
  assign regs_io_argOuts_54_bits = {{32'd0}, mags_0_io_debugSignals_52};
  assign regs_io_argOuts_55_bits = {{32'd0}, mags_0_io_debugSignals_53};
  assign regs_io_argOuts_56_bits = {{32'd0}, mags_0_io_debugSignals_54};
  assign regs_io_argOuts_57_bits = {{32'd0}, mags_0_io_debugSignals_55};
  assign regs_io_argOuts_58_bits = {{32'd0}, mags_0_io_debugSignals_56};
  assign regs_io_argOuts_59_bits = {{32'd0}, mags_0_io_debugSignals_57};
  assign regs_io_argOuts_60_bits = {{32'd0}, mags_0_io_debugSignals_58};
  assign regs_clock = clock;
  assign regs_reset = reset;
  assign timeoutCtr_io_max = 40'h2cb417800;
  assign timeoutCtr_io_enable = localEnable;
  assign timeoutCtr_io_saturate = 1'h1;
  assign timeoutCtr_clock = clock;
  assign timeoutCtr_reset = reset;
  assign depulser_io_in = _T_358;
  assign depulser_io_rst = _T_359[0];
  assign depulser_clock = clock;
  assign depulser_reset = reset;
  assign status_valid = depulser_io_out;
  assign status_bits = {{62'd0}, _T_372};
endmodule
module FringeArria10(
  input         clock,
  input         reset,
  output [31:0] io_S_AVALON_readdata,
  input  [7:0]  io_S_AVALON_address,
  input         io_S_AVALON_write,
  input  [31:0] io_S_AVALON_writedata,
  output        io_enable,
  input         io_done,
  output [31:0] io_argIns_0,
  input         io_argOuts_0_valid,
  input  [31:0] io_argOuts_0_bits
);
  wire  fringeCommon_clock;
  wire  fringeCommon_reset;
  wire [31:0] fringeCommon_io_raddr;
  wire  fringeCommon_io_wen;
  wire [31:0] fringeCommon_io_waddr;
  wire [63:0] fringeCommon_io_wdata;
  wire [63:0] fringeCommon_io_rdata;
  wire  fringeCommon_io_enable;
  wire  fringeCommon_io_done;
  wire [63:0] fringeCommon_io_argIns_0;
  wire  fringeCommon_io_argOuts_0_valid;
  wire [63:0] fringeCommon_io_argOuts_0_bits;
  Fringe fringeCommon (
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits)
  );
  assign io_S_AVALON_readdata = fringeCommon_io_rdata[31:0];
  assign io_enable = fringeCommon_io_enable;
  assign io_argIns_0 = fringeCommon_io_argIns_0[31:0];
  assign fringeCommon_io_raddr = {{24'd0}, io_S_AVALON_address};
  assign fringeCommon_io_wen = io_S_AVALON_write;
  assign fringeCommon_io_waddr = {{24'd0}, io_S_AVALON_address};
  assign fringeCommon_io_wdata = {{32'd0}, io_S_AVALON_writedata};
  assign fringeCommon_io_done = io_done;
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid;
  assign fringeCommon_io_argOuts_0_bits = {{32'd0}, io_argOuts_0_bits};
  assign fringeCommon_clock = clock;
  assign fringeCommon_reset = reset;
endmodule
module Top(
  input         clock,
  input         reset,
  input         io_raddr,
  input         io_wen,
  input         io_waddr,
  input         io_wdata,
  output        io_rdata,
  output [31:0] io_S_AVALON_readdata,
  input  [7:0]  io_S_AVALON_address,
  input         io_S_AVALON_chipselect,
  input         io_S_AVALON_write,
  input         io_S_AVALON_read,
  input  [31:0] io_S_AVALON_writedata
);
  wire  accel_clock;
  wire  accel_reset;
  wire  accel_io_enable;
  wire  accel_io_done;
  wire [63:0] accel_io_argIns_0;
  wire  accel_io_argOuts_0_valid;
  wire [63:0] accel_io_argOuts_0_bits;
  wire  FringeArria10_clock;
  wire  FringeArria10_reset;
  wire [31:0] FringeArria10_io_S_AVALON_readdata;
  wire [7:0] FringeArria10_io_S_AVALON_address;
  wire  FringeArria10_io_S_AVALON_write;
  wire [31:0] FringeArria10_io_S_AVALON_writedata;
  wire  FringeArria10_io_enable;
  wire  FringeArria10_io_done;
  wire [31:0] FringeArria10_io_argIns_0;
  wire  FringeArria10_io_argOuts_0_valid;
  wire [31:0] FringeArria10_io_argOuts_0_bits;
  AccelTop accel (
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_argIns_0(accel_io_argIns_0),
    .io_argOuts_0_valid(accel_io_argOuts_0_valid),
    .io_argOuts_0_bits(accel_io_argOuts_0_bits)
  );
  FringeArria10 FringeArria10 (
    .clock(FringeArria10_clock),
    .reset(FringeArria10_reset),
    .io_S_AVALON_readdata(FringeArria10_io_S_AVALON_readdata),
    .io_S_AVALON_address(FringeArria10_io_S_AVALON_address),
    .io_S_AVALON_write(FringeArria10_io_S_AVALON_write),
    .io_S_AVALON_writedata(FringeArria10_io_S_AVALON_writedata),
    .io_enable(FringeArria10_io_enable),
    .io_done(FringeArria10_io_done),
    .io_argIns_0(FringeArria10_io_argIns_0),
    .io_argOuts_0_valid(FringeArria10_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeArria10_io_argOuts_0_bits)
  );
  assign io_rdata = 1'h0;
  assign io_S_AVALON_readdata = FringeArria10_io_S_AVALON_readdata;
  assign accel_io_enable = FringeArria10_io_enable;
  assign accel_io_argIns_0 = {{32'd0}, FringeArria10_io_argIns_0};
  assign accel_clock = clock;
  assign accel_reset = reset;
  assign FringeArria10_io_S_AVALON_address = io_S_AVALON_address;
  assign FringeArria10_io_S_AVALON_write = io_S_AVALON_write;
  assign FringeArria10_io_S_AVALON_writedata = io_S_AVALON_writedata;
  assign FringeArria10_io_done = accel_io_done;
  assign FringeArria10_io_argOuts_0_valid = accel_io_argOuts_0_valid;
  assign FringeArria10_io_argOuts_0_bits = accel_io_argOuts_0_bits[31:0];
  assign FringeArria10_clock = clock;
  assign FringeArria10_reset = reset;
endmodule
